`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/29/2025 09:15:25 PM
// Design Name: 
// Module Name: game_over
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module game_over
	(
		input clk,
		input [9:0] row,
		input [9:0] col,
		output reg [11:0] color_data,
		input ce
	);
	    (* rom_style = "block" *)
	    
	reg [9:0] row_reg;
	reg [9:0] col_reg;
	always @(posedge clk)
		begin
		if (ce) begin
		row_reg <= row;
		col_reg <= col;
		end
		end
	always @(*) begin
	case ({row_reg, col_reg})
		20'b00101001010011110010: color_data = 12'b000000010000;
20'b00101001010011110011: color_data = 12'b000000010000;
20'b00101001010011110100: color_data = 12'b000000010000;
20'b00101001010100101000: color_data = 12'b000000000010;
20'b00101001010100101001: color_data = 12'b000000000011;
20'b00101001010100101010: color_data = 12'b000000000011;
20'b00101001010100101011: color_data = 12'b000000000010;
20'b00101001010100101100: color_data = 12'b000000000010;
20'b00101001010100101101: color_data = 12'b000000000010;
20'b00101001010100101110: color_data = 12'b000000000010;
20'b00101001010100101111: color_data = 12'b000000000010;
20'b00101001010100110000: color_data = 12'b000000000010;
20'b00101001010100110001: color_data = 12'b000000000010;
20'b00101001100011110000: color_data = 12'b000000010000;
20'b00101001100011110001: color_data = 12'b011011011010;
20'b00101001100011110010: color_data = 12'b001111101001;
20'b00101001100011110011: color_data = 12'b001111111001;
20'b00101001100011110100: color_data = 12'b001111101001;
20'b00101001100011110101: color_data = 12'b010111101010;
20'b00101001100011110110: color_data = 12'b000000010000;
20'b00101001100100100111: color_data = 12'b000000000010;
20'b00101001100100101000: color_data = 12'b001000011011;
20'b00101001100100101001: color_data = 12'b000100011101;
20'b00101001100100101010: color_data = 12'b000000001100;
20'b00101001100100101011: color_data = 12'b000100011100;
20'b00101001100100101100: color_data = 12'b000000000101;
20'b00101001100100101101: color_data = 12'b001000101010;
20'b00101001100100101110: color_data = 12'b000100011011;
20'b00101001100100101111: color_data = 12'b000100011101;
20'b00101001100100110000: color_data = 12'b000100011100;
20'b00101001100100110001: color_data = 12'b000100011010;
20'b00101001100100110010: color_data = 12'b000000000010;
20'b00101001110011110000: color_data = 12'b000000010000;
20'b00101001110011110001: color_data = 12'b010011101001;
20'b00101001110011110010: color_data = 12'b000111111000;
20'b00101001110011110011: color_data = 12'b000011111000;
20'b00101001110011110100: color_data = 12'b000011111000;
20'b00101001110011110101: color_data = 12'b001111101001;
20'b00101001110011110110: color_data = 12'b000000010000;
20'b00101001110100100111: color_data = 12'b000000000010;
20'b00101001110100101000: color_data = 12'b000100011101;
20'b00101001110100101001: color_data = 12'b000000001111;
20'b00101001110100101010: color_data = 12'b000000001111;
20'b00101001110100101011: color_data = 12'b000000001110;
20'b00101001110100101100: color_data = 12'b000000000110;
20'b00101001110100101101: color_data = 12'b000100011011;
20'b00101001110100101110: color_data = 12'b000100001110;
20'b00101001110100101111: color_data = 12'b000000001111;
20'b00101001110100110000: color_data = 12'b000000001111;
20'b00101001110100110001: color_data = 12'b000100011100;
20'b00101001110100110010: color_data = 12'b000000000010;
20'b00101001110101110000: color_data = 12'b000000010000;
20'b00101001110101110001: color_data = 12'b000000010000;
20'b00101001110101110010: color_data = 12'b000000010000;
20'b00101001110101111000: color_data = 12'b000000010000;
20'b00101010000011110000: color_data = 12'b000000010000;
20'b00101010000011110001: color_data = 12'b010011101001;
20'b00101010000011110010: color_data = 12'b000111111000;
20'b00101010000011110011: color_data = 12'b000011111000;
20'b00101010000011110100: color_data = 12'b000011110111;
20'b00101010000011110101: color_data = 12'b001111111000;
20'b00101010000011110110: color_data = 12'b000000010000;
20'b00101010000100100111: color_data = 12'b000000000010;
20'b00101010000100101000: color_data = 12'b000100011101;
20'b00101010000100101001: color_data = 12'b000000001111;
20'b00101010000100101010: color_data = 12'b000000001111;
20'b00101010000100101011: color_data = 12'b000000001110;
20'b00101010000100101100: color_data = 12'b000000000110;
20'b00101010000100101101: color_data = 12'b000100101011;
20'b00101010000100101110: color_data = 12'b000000001110;
20'b00101010000100101111: color_data = 12'b000000001111;
20'b00101010000100110000: color_data = 12'b000000001111;
20'b00101010000100110001: color_data = 12'b000000011100;
20'b00101010000100110010: color_data = 12'b000000000010;
20'b00101010000101101111: color_data = 12'b011011011010;
20'b00101010000101110000: color_data = 12'b001111101001;
20'b00101010000101110001: color_data = 12'b001011101000;
20'b00101010000101110010: color_data = 12'b001011101001;
20'b00101010000101110011: color_data = 12'b010011101001;
20'b00101010000101110100: color_data = 12'b000000100000;
20'b00101010000101110101: color_data = 12'b011011011010;
20'b00101010000101110110: color_data = 12'b010011101001;
20'b00101010000101110111: color_data = 12'b001111101001;
20'b00101010000101111000: color_data = 12'b001011101001;
20'b00101010000101111001: color_data = 12'b010111101001;
20'b00101010000101111010: color_data = 12'b000000010000;
20'b00101010010011101111: color_data = 12'b000000010000;
20'b00101010010011110000: color_data = 12'b000000010000;
20'b00101010010011110001: color_data = 12'b010111101001;
20'b00101010010011110010: color_data = 12'b001011111000;
20'b00101010010011110011: color_data = 12'b000011110111;
20'b00101010010011110100: color_data = 12'b000111111000;
20'b00101010010011110101: color_data = 12'b010011101001;
20'b00101010010011110110: color_data = 12'b000000010000;
20'b00101010010100100111: color_data = 12'b000000000010;
20'b00101010010100101000: color_data = 12'b001000011010;
20'b00101010010100101001: color_data = 12'b000100011100;
20'b00101010010100101010: color_data = 12'b000100011100;
20'b00101010010100101011: color_data = 12'b000100011011;
20'b00101010010100101100: color_data = 12'b000000000101;
20'b00101010010100101101: color_data = 12'b000100101010;
20'b00101010010100101110: color_data = 12'b000000011101;
20'b00101010010100101111: color_data = 12'b000000001110;
20'b00101010010100110000: color_data = 12'b000000001110;
20'b00101010010100110001: color_data = 12'b000100011011;
20'b00101010010100110010: color_data = 12'b000000000010;
20'b00101010010101101110: color_data = 12'b000000010000;
20'b00101010010101101111: color_data = 12'b010011011010;
20'b00101010010101110000: color_data = 12'b000011111000;
20'b00101010010101110001: color_data = 12'b000011111000;
20'b00101010010101110010: color_data = 12'b000011110111;
20'b00101010010101110011: color_data = 12'b000111111000;
20'b00101010010101110100: color_data = 12'b000000100000;
20'b00101010010101110101: color_data = 12'b010011101001;
20'b00101010010101110110: color_data = 12'b001011111000;
20'b00101010010101110111: color_data = 12'b000011110111;
20'b00101010010101111000: color_data = 12'b000011111000;
20'b00101010010101111001: color_data = 12'b001011101000;
20'b00101010010101111010: color_data = 12'b000000010000;
20'b00101010100011101011: color_data = 12'b000000010000;
20'b00101010100011101100: color_data = 12'b000000010000;
20'b00101010100011101101: color_data = 12'b000000010000;
20'b00101010100011101110: color_data = 12'b000000100000;
20'b00101010100011101111: color_data = 12'b000000010000;
20'b00101010100011110000: color_data = 12'b000000010000;
20'b00101010100011110001: color_data = 12'b000000010000;
20'b00101010100011110010: color_data = 12'b000000100000;
20'b00101010100011110011: color_data = 12'b000000100000;
20'b00101010100011110100: color_data = 12'b000000110000;
20'b00101010100011110101: color_data = 12'b000000100000;
20'b00101010100100101000: color_data = 12'b000000000010;
20'b00101010100100101001: color_data = 12'b000000000010;
20'b00101010100100101010: color_data = 12'b000000000011;
20'b00101010100100101011: color_data = 12'b000000000010;
20'b00101010100100101100: color_data = 12'b000000000011;
20'b00101010100100101101: color_data = 12'b000000000100;
20'b00101010100100101110: color_data = 12'b000000000101;
20'b00101010100100101111: color_data = 12'b000000000111;
20'b00101010100100110000: color_data = 12'b000000000111;
20'b00101010100100110001: color_data = 12'b000000000101;
20'b00101010100100110010: color_data = 12'b000000000001;
20'b00101010100101101110: color_data = 12'b000000010000;
20'b00101010100101101111: color_data = 12'b010011101010;
20'b00101010100101110000: color_data = 12'b000111111000;
20'b00101010100101110001: color_data = 12'b000011110111;
20'b00101010100101110010: color_data = 12'b000011110111;
20'b00101010100101110011: color_data = 12'b000111111000;
20'b00101010100101110100: color_data = 12'b000000100000;
20'b00101010100101110101: color_data = 12'b010011101001;
20'b00101010100101110110: color_data = 12'b000111111000;
20'b00101010100101110111: color_data = 12'b000011111000;
20'b00101010100101111000: color_data = 12'b000011110111;
20'b00101010100101111001: color_data = 12'b001111111001;
20'b00101010100101111010: color_data = 12'b000000010000;
20'b00101010110011101001: color_data = 12'b000000010000;
20'b00101010110011101010: color_data = 12'b000000010000;
20'b00101010110011101011: color_data = 12'b011111011010;
20'b00101010110011101100: color_data = 12'b010111101010;
20'b00101010110011101101: color_data = 12'b010011011001;
20'b00101010110011101110: color_data = 12'b010011101001;
20'b00101010110011101111: color_data = 12'b010111101001;
20'b00101010110011110000: color_data = 12'b000000010000;
20'b00101010110011110001: color_data = 12'b011111011001;
20'b00101010110011110010: color_data = 12'b010111101001;
20'b00101010110011110011: color_data = 12'b010011101001;
20'b00101010110011110100: color_data = 12'b001111101001;
20'b00101010110011110101: color_data = 12'b010111011010;
20'b00101010110011110110: color_data = 12'b000000010000;
20'b00101010110100101011: color_data = 12'b000000000001;
20'b00101010110100101100: color_data = 12'b000000000010;
20'b00101010110100101101: color_data = 12'b001100111001;
20'b00101010110100101110: color_data = 12'b001000101010;
20'b00101010110100101111: color_data = 12'b000100011011;
20'b00101010110100110000: color_data = 12'b001000011011;
20'b00101010110100110001: color_data = 12'b001000101001;
20'b00101010110100110010: color_data = 12'b000000000001;
20'b00101010110101101110: color_data = 12'b000000010000;
20'b00101010110101101111: color_data = 12'b010111101010;
20'b00101010110101110000: color_data = 12'b001111111001;
20'b00101010110101110001: color_data = 12'b000111111000;
20'b00101010110101110010: color_data = 12'b000111111000;
20'b00101010110101110011: color_data = 12'b001111111000;
20'b00101010110101110100: color_data = 12'b000000100000;
20'b00101010110101110101: color_data = 12'b010111101001;
20'b00101010110101110110: color_data = 12'b001011101000;
20'b00101010110101110111: color_data = 12'b000111111000;
20'b00101010110101111000: color_data = 12'b000111111000;
20'b00101010110101111001: color_data = 12'b010011101000;
20'b00101011000011101010: color_data = 12'b000000010000;
20'b00101011000011101011: color_data = 12'b010111011001;
20'b00101011000011101100: color_data = 12'b001111101001;
20'b00101011000011101101: color_data = 12'b001011111001;
20'b00101011000011101110: color_data = 12'b000111111000;
20'b00101011000011101111: color_data = 12'b001011101000;
20'b00101011000011110000: color_data = 12'b000000100000;
20'b00101011000011110001: color_data = 12'b010111101001;
20'b00101011000011110010: color_data = 12'b001011101000;
20'b00101011000011110011: color_data = 12'b000111111000;
20'b00101011000011110100: color_data = 12'b000011111000;
20'b00101011000011110101: color_data = 12'b001111101001;
20'b00101011000100101011: color_data = 12'b000000000001;
20'b00101011000100101100: color_data = 12'b000000000011;
20'b00101011000100101101: color_data = 12'b001000101011;
20'b00101011000100101110: color_data = 12'b000100011101;
20'b00101011000100101111: color_data = 12'b000100001110;
20'b00101011000100110000: color_data = 12'b000000001110;
20'b00101011000100110001: color_data = 12'b001000011100;
20'b00101011000100110010: color_data = 12'b000000000010;
20'b00101011000101101110: color_data = 12'b000000010000;
20'b00101011000101101111: color_data = 12'b011011011001;
20'b00101011000101110000: color_data = 12'b010111011001;
20'b00101011000101110001: color_data = 12'b010011011000;
20'b00101011000101110010: color_data = 12'b010011101001;
20'b00101011000101110011: color_data = 12'b010111101001;
20'b00101011000101110100: color_data = 12'b000000010000;
20'b00101011000101110101: color_data = 12'b011111011010;
20'b00101011000101110110: color_data = 12'b010011011010;
20'b00101011000101110111: color_data = 12'b001111101001;
20'b00101011000101111000: color_data = 12'b010011101001;
20'b00101011000101111001: color_data = 12'b011011101010;
20'b00101011010011101001: color_data = 12'b000000010000;
20'b00101011010011101010: color_data = 12'b000000010000;
20'b00101011010011101011: color_data = 12'b010011101001;
20'b00101011010011101100: color_data = 12'b000111111001;
20'b00101011010011101101: color_data = 12'b000011111000;
20'b00101011010011101110: color_data = 12'b000011111000;
20'b00101011010011101111: color_data = 12'b000111111000;
20'b00101011010011110000: color_data = 12'b000000100000;
20'b00101011010011110001: color_data = 12'b010011101001;
20'b00101011010011110010: color_data = 12'b000111111000;
20'b00101011010011110011: color_data = 12'b000011111000;
20'b00101011010011110100: color_data = 12'b000011111000;
20'b00101011010011110101: color_data = 12'b001111111001;
20'b00101011010011110110: color_data = 12'b000000010000;
20'b00101011010100101011: color_data = 12'b000000000001;
20'b00101011010100101100: color_data = 12'b000000000100;
20'b00101011010100101101: color_data = 12'b001000011011;
20'b00101011010100101110: color_data = 12'b000000001110;
20'b00101011010100101111: color_data = 12'b000000001111;
20'b00101011010100110000: color_data = 12'b000000001111;
20'b00101011010100110001: color_data = 12'b000100011101;
20'b00101011010100110010: color_data = 12'b000000000011;
20'b00101011010101101110: color_data = 12'b000000010000;
20'b00101011010101101111: color_data = 12'b000000010000;
20'b00101011010101110000: color_data = 12'b000000100000;
20'b00101011010101110001: color_data = 12'b000000100000;
20'b00101011010101110010: color_data = 12'b000000100000;
20'b00101011010101110011: color_data = 12'b000000100000;
20'b00101011010101110100: color_data = 12'b000000010000;
20'b00101011010101110110: color_data = 12'b000000010000;
20'b00101011010101110111: color_data = 12'b000000010000;
20'b00101011010101111000: color_data = 12'b000000010000;
20'b00101011010101111001: color_data = 12'b000000010000;
20'b00101011100011101010: color_data = 12'b000000010000;
20'b00101011100011101011: color_data = 12'b010011101001;
20'b00101011100011101100: color_data = 12'b000111111000;
20'b00101011100011101101: color_data = 12'b000011111000;
20'b00101011100011101110: color_data = 12'b000011110111;
20'b00101011100011101111: color_data = 12'b000111111000;
20'b00101011100011110000: color_data = 12'b000000100000;
20'b00101011100011110001: color_data = 12'b010011101001;
20'b00101011100011110010: color_data = 12'b000111111000;
20'b00101011100011110011: color_data = 12'b000011111000;
20'b00101011100011110100: color_data = 12'b000011110111;
20'b00101011100011110101: color_data = 12'b001011101000;
20'b00101011100011110110: color_data = 12'b000000010000;
20'b00101011100100101011: color_data = 12'b000000000001;
20'b00101011100100101100: color_data = 12'b000000000100;
20'b00101011100100101101: color_data = 12'b000100011100;
20'b00101011100100101110: color_data = 12'b000000001110;
20'b00101011100100101111: color_data = 12'b000000001111;
20'b00101011100100110000: color_data = 12'b000000001111;
20'b00101011100100110001: color_data = 12'b000100011101;
20'b00101011100100110010: color_data = 12'b000000000010;
20'b00101011100101101110: color_data = 12'b000000010000;
20'b00101011100101101111: color_data = 12'b010111101001;
20'b00101011100101110000: color_data = 12'b001011101000;
20'b00101011100101110001: color_data = 12'b000111111000;
20'b00101011100101110010: color_data = 12'b000111111000;
20'b00101011100101110011: color_data = 12'b010011101001;
20'b00101011100101110100: color_data = 12'b000000010000;
20'b00101011110011101010: color_data = 12'b000000010000;
20'b00101011110011101011: color_data = 12'b011011011010;
20'b00101011110011101100: color_data = 12'b001111101001;
20'b00101011110011101101: color_data = 12'b001011101001;
20'b00101011110011101110: color_data = 12'b001111111000;
20'b00101011110011101111: color_data = 12'b010011101001;
20'b00101011110011110000: color_data = 12'b000000010000;
20'b00101011110011110001: color_data = 12'b011011101010;
20'b00101011110011110010: color_data = 12'b001111101001;
20'b00101011110011110011: color_data = 12'b001011101000;
20'b00101011110011110100: color_data = 12'b001011111001;
20'b00101011110011110101: color_data = 12'b010011101001;
20'b00101011110011110110: color_data = 12'b000000010000;
20'b00101011110100101011: color_data = 12'b000000000001;
20'b00101011110100101100: color_data = 12'b000000000011;
20'b00101011110100101101: color_data = 12'b001000101010;
20'b00101011110100101110: color_data = 12'b000100011011;
20'b00101011110100101111: color_data = 12'b000000011100;
20'b00101011110100110000: color_data = 12'b000000011100;
20'b00101011110100110001: color_data = 12'b000100101010;
20'b00101011110100110010: color_data = 12'b000000000010;
20'b00101011110101000100: color_data = 12'b000100000000;
20'b00101011110101000101: color_data = 12'b000100000000;
20'b00101011110101000110: color_data = 12'b000100000000;
20'b00101011110101000111: color_data = 12'b000100000000;
20'b00101011110101001000: color_data = 12'b000100000000;
20'b00101011110101001001: color_data = 12'b000100000000;
20'b00101011110101001010: color_data = 12'b000100000000;
20'b00101011110101001011: color_data = 12'b000100000000;
20'b00101011110101001100: color_data = 12'b000100000000;
20'b00101011110101001101: color_data = 12'b000100000000;
20'b00101011110101101110: color_data = 12'b000000010000;
20'b00101011110101101111: color_data = 12'b010011101001;
20'b00101011110101110000: color_data = 12'b000111111000;
20'b00101011110101110001: color_data = 12'b000011111000;
20'b00101011110101110010: color_data = 12'b000011110111;
20'b00101011110101110011: color_data = 12'b001111111000;
20'b00101011110101110100: color_data = 12'b000000010000;
20'b00101100000011101101: color_data = 12'b000000010000;
20'b00101100000011101110: color_data = 12'b000000010000;
20'b00101100000011110011: color_data = 12'b000000010000;
20'b00101100000011110100: color_data = 12'b000000010000;
20'b00101100000100101100: color_data = 12'b000000000001;
20'b00101100000100101101: color_data = 12'b000000000001;
20'b00101100000100101110: color_data = 12'b000000000010;
20'b00101100000100101111: color_data = 12'b000000000010;
20'b00101100000100110000: color_data = 12'b000000000010;
20'b00101100000100110001: color_data = 12'b000000000001;
20'b00101100000101000010: color_data = 12'b000100000000;
20'b00101100000101000011: color_data = 12'b001000000000;
20'b00101100000101000100: color_data = 12'b010000000000;
20'b00101100000101000101: color_data = 12'b010100000000;
20'b00101100000101000110: color_data = 12'b010100000000;
20'b00101100000101000111: color_data = 12'b010000000000;
20'b00101100000101001000: color_data = 12'b001100000000;
20'b00101100000101001001: color_data = 12'b001100000000;
20'b00101100000101001010: color_data = 12'b010000000000;
20'b00101100000101001011: color_data = 12'b010100000000;
20'b00101100000101001100: color_data = 12'b010100000000;
20'b00101100000101001101: color_data = 12'b001100000000;
20'b00101100000101001110: color_data = 12'b000100000000;
20'b00101100000101101110: color_data = 12'b000000010000;
20'b00101100000101101111: color_data = 12'b010011101001;
20'b00101100000101110000: color_data = 12'b000111111000;
20'b00101100000101110001: color_data = 12'b000011110111;
20'b00101100000101110010: color_data = 12'b000011110111;
20'b00101100000101110011: color_data = 12'b001011111000;
20'b00101100000101110100: color_data = 12'b000000010000;
20'b00101100010101000010: color_data = 12'b001000000000;
20'b00101100010101000011: color_data = 12'b011000010000;
20'b00101100010101000100: color_data = 12'b100100000000;
20'b00101100010101000101: color_data = 12'b101000000000;
20'b00101100010101000110: color_data = 12'b101000000000;
20'b00101100010101000111: color_data = 12'b100100000000;
20'b00101100010101001000: color_data = 12'b010100000000;
20'b00101100010101001001: color_data = 12'b011100010001;
20'b00101100010101001010: color_data = 12'b100100000000;
20'b00101100010101001011: color_data = 12'b101000000000;
20'b00101100010101001100: color_data = 12'b101000000000;
20'b00101100010101001101: color_data = 12'b100000000000;
20'b00101100010101001110: color_data = 12'b001000000000;
20'b00101100010101101110: color_data = 12'b000000010000;
20'b00101100010101101111: color_data = 12'b010111101010;
20'b00101100010101110000: color_data = 12'b001011101001;
20'b00101100010101110001: color_data = 12'b000111111000;
20'b00101100010101110010: color_data = 12'b000111111000;
20'b00101100010101110011: color_data = 12'b001111101000;
20'b00101100010101110100: color_data = 12'b000000010000;
20'b00101100100101000001: color_data = 12'b000100000000;
20'b00101100100101000010: color_data = 12'b010000000000;
20'b00101100100101000011: color_data = 12'b100100010000;
20'b00101100100101000100: color_data = 12'b110000000000;
20'b00101100100101000101: color_data = 12'b111000000000;
20'b00101100100101000110: color_data = 12'b111000000000;
20'b00101100100101000111: color_data = 12'b110000000000;
20'b00101100100101001000: color_data = 12'b011100000000;
20'b00101100100101001001: color_data = 12'b100100000000;
20'b00101100100101001010: color_data = 12'b110000000000;
20'b00101100100101001011: color_data = 12'b111000000000;
20'b00101100100101001100: color_data = 12'b110100000000;
20'b00101100100101001101: color_data = 12'b101100000000;
20'b00101100100101001110: color_data = 12'b001100000000;
20'b00101100100101101110: color_data = 12'b000000010000;
20'b00101100100101101111: color_data = 12'b000000010000;
20'b00101100100101110000: color_data = 12'b000000100000;
20'b00101100100101110001: color_data = 12'b000000100000;
20'b00101100100101110010: color_data = 12'b000000100000;
20'b00101100100101110011: color_data = 12'b000000100000;
20'b00101100110101000001: color_data = 12'b000100000000;
20'b00101100110101000010: color_data = 12'b010000000000;
20'b00101100110101000011: color_data = 12'b100100000000;
20'b00101100110101000100: color_data = 12'b110000000000;
20'b00101100110101000101: color_data = 12'b111000000000;
20'b00101100110101000110: color_data = 12'b110100000000;
20'b00101100110101000111: color_data = 12'b110000000000;
20'b00101100110101001000: color_data = 12'b011100000000;
20'b00101100110101001001: color_data = 12'b100100010001;
20'b00101100110101001010: color_data = 12'b110000000000;
20'b00101100110101001011: color_data = 12'b110100000000;
20'b00101100110101001100: color_data = 12'b110100000000;
20'b00101100110101001101: color_data = 12'b101100000000;
20'b00101100110101001110: color_data = 12'b001100000000;
20'b00101100110101101110: color_data = 12'b000000010000;
20'b00101100110101101111: color_data = 12'b011111011010;
20'b00101100110101110000: color_data = 12'b010111011001;
20'b00101100110101110001: color_data = 12'b010011101001;
20'b00101100110101110010: color_data = 12'b010011101001;
20'b00101100110101110011: color_data = 12'b011011011010;
20'b00101101000101000001: color_data = 12'b000100000000;
20'b00101101000101000010: color_data = 12'b001100000000;
20'b00101101000101000011: color_data = 12'b011100010001;
20'b00101101000101000100: color_data = 12'b100100000000;
20'b00101101000101000101: color_data = 12'b101000000000;
20'b00101101000101000110: color_data = 12'b101000000000;
20'b00101101000101000111: color_data = 12'b100100000001;
20'b00101101000101001000: color_data = 12'b010100000000;
20'b00101101000101001001: color_data = 12'b011100000000;
20'b00101101000101001010: color_data = 12'b101000010000;
20'b00101101000101001011: color_data = 12'b101000000000;
20'b00101101000101001100: color_data = 12'b101000010000;
20'b00101101000101001101: color_data = 12'b100000010000;
20'b00101101000101001110: color_data = 12'b001000000000;
20'b00101101000101101110: color_data = 12'b000000010000;
20'b00101101000101101111: color_data = 12'b010111011001;
20'b00101101000101110000: color_data = 12'b001011111001;
20'b00101101000101110001: color_data = 12'b000111111000;
20'b00101101000101110010: color_data = 12'b001011111000;
20'b00101101000101110011: color_data = 12'b010011101001;
20'b00101101000101110100: color_data = 12'b000000010000;
20'b00101101010101000001: color_data = 12'b000100000000;
20'b00101101010101000010: color_data = 12'b001000000000;
20'b00101101010101000011: color_data = 12'b001100000000;
20'b00101101010101000100: color_data = 12'b010000000000;
20'b00101101010101000101: color_data = 12'b010100000000;
20'b00101101010101000110: color_data = 12'b010100000000;
20'b00101101010101000111: color_data = 12'b010100000000;
20'b00101101010101001000: color_data = 12'b010000000000;
20'b00101101010101001001: color_data = 12'b010100000000;
20'b00101101010101001010: color_data = 12'b100000000000;
20'b00101101010101001011: color_data = 12'b100000000000;
20'b00101101010101001100: color_data = 12'b100000000000;
20'b00101101010101001101: color_data = 12'b011000000000;
20'b00101101010101001110: color_data = 12'b001100000000;
20'b00101101010101001111: color_data = 12'b001000000000;
20'b00101101010101010000: color_data = 12'b001100000000;
20'b00101101010101010001: color_data = 12'b001100000000;
20'b00101101010101010010: color_data = 12'b001000000000;
20'b00101101010101010011: color_data = 12'b000100000000;
20'b00101101010101101110: color_data = 12'b000000010000;
20'b00101101010101101111: color_data = 12'b010111011010;
20'b00101101010101110000: color_data = 12'b001011101001;
20'b00101101010101110001: color_data = 12'b000111111000;
20'b00101101010101110010: color_data = 12'b000111111000;
20'b00101101010101110011: color_data = 12'b010011101001;
20'b00101101010101110100: color_data = 12'b000000010000;
20'b00101101100011110110: color_data = 12'b111111111111;
20'b00101101100011110111: color_data = 12'b111011101110;
20'b00101101100011111000: color_data = 12'b111011101110;
20'b00101101100011111001: color_data = 12'b111011101110;
20'b00101101100011111010: color_data = 12'b111111111111;
20'b00101101100011111100: color_data = 12'b111011101110;
20'b00101101100011111101: color_data = 12'b111011101110;
20'b00101101100011111110: color_data = 12'b111011101110;
20'b00101101100011111111: color_data = 12'b111011101110;
20'b00101101100100000001: color_data = 12'b111011101110;
20'b00101101100100000010: color_data = 12'b111111111111;
20'b00101101100100000011: color_data = 12'b111011101110;
20'b00101101100100000100: color_data = 12'b111011101110;
20'b00101101100100000101: color_data = 12'b111111111111;
20'b00101101100100000111: color_data = 12'b111011101110;
20'b00101101100100001000: color_data = 12'b111011101110;
20'b00101101100100001001: color_data = 12'b111011101110;
20'b00101101100100001010: color_data = 12'b111011101110;
20'b00101101100100001011: color_data = 12'b111011101110;
20'b00101101100100100011: color_data = 12'b111011101110;
20'b00101101100100100100: color_data = 12'b111111111111;
20'b00101101100100100101: color_data = 12'b111011101110;
20'b00101101100100100110: color_data = 12'b111011101110;
20'b00101101100101000011: color_data = 12'b000100000000;
20'b00101101100101000100: color_data = 12'b000100000000;
20'b00101101100101000101: color_data = 12'b000100000000;
20'b00101101100101000110: color_data = 12'b000100000000;
20'b00101101100101000111: color_data = 12'b001000000000;
20'b00101101100101001000: color_data = 12'b010100000000;
20'b00101101100101001001: color_data = 12'b100100000000;
20'b00101101100101001010: color_data = 12'b110000000000;
20'b00101101100101001011: color_data = 12'b110100000000;
20'b00101101100101001100: color_data = 12'b111000000000;
20'b00101101100101001101: color_data = 12'b110000000000;
20'b00101101100101001110: color_data = 12'b011100000000;
20'b00101101100101001111: color_data = 12'b100000000001;
20'b00101101100101010000: color_data = 12'b101100000000;
20'b00101101100101010001: color_data = 12'b101000000000;
20'b00101101100101010010: color_data = 12'b100000000000;
20'b00101101100101010011: color_data = 12'b010000000000;
20'b00101101100101010100: color_data = 12'b000100000000;
20'b00101101100101011111: color_data = 12'b111011101110;
20'b00101101100101100000: color_data = 12'b111111101110;
20'b00101101100101100001: color_data = 12'b111011101110;
20'b00101101100101100010: color_data = 12'b111111111111;
20'b00101101100101100100: color_data = 12'b111011101110;
20'b00101101100101100101: color_data = 12'b111111101110;
20'b00101101100101100110: color_data = 12'b111011101110;
20'b00101101100101100111: color_data = 12'b111111101110;
20'b00101101100101101000: color_data = 12'b111011101110;
20'b00101101100101101111: color_data = 12'b011111011010;
20'b00101101100101110000: color_data = 12'b010111101001;
20'b00101101100101110001: color_data = 12'b010011101001;
20'b00101101100101110010: color_data = 12'b010011101001;
20'b00101101100101110011: color_data = 12'b011111101001;
20'b00101101110011110110: color_data = 12'b111011101110;
20'b00101101110011110111: color_data = 12'b111011101110;
20'b00101101110011111000: color_data = 12'b111011101110;
20'b00101101110011111001: color_data = 12'b111111111111;
20'b00101101110011111010: color_data = 12'b111011101110;
20'b00101101110011111100: color_data = 12'b111011101110;
20'b00101101110011111101: color_data = 12'b111011101110;
20'b00101101110011111110: color_data = 12'b111011101110;
20'b00101101110011111111: color_data = 12'b111011101110;
20'b00101101110100000001: color_data = 12'b111011101110;
20'b00101101110100000010: color_data = 12'b111111111111;
20'b00101101110100000011: color_data = 12'b111011101110;
20'b00101101110100000100: color_data = 12'b111011101110;
20'b00101101110100000101: color_data = 12'b111011101110;
20'b00101101110100000111: color_data = 12'b111011101110;
20'b00101101110100001000: color_data = 12'b111011101110;
20'b00101101110100001001: color_data = 12'b111011101110;
20'b00101101110100001010: color_data = 12'b111011101110;
20'b00101101110100001011: color_data = 12'b111011101110;
20'b00101101110100100011: color_data = 12'b111011101110;
20'b00101101110100100100: color_data = 12'b111011101110;
20'b00101101110100100101: color_data = 12'b111011101110;
20'b00101101110100100110: color_data = 12'b111011101110;
20'b00101101110101000111: color_data = 12'b000100000000;
20'b00101101110101001000: color_data = 12'b010100000000;
20'b00101101110101001001: color_data = 12'b101000000000;
20'b00101101110101001010: color_data = 12'b110100000000;
20'b00101101110101001011: color_data = 12'b111100000000;
20'b00101101110101001100: color_data = 12'b111100000000;
20'b00101101110101001101: color_data = 12'b110100000000;
20'b00101101110101001110: color_data = 12'b100100000000;
20'b00101101110101001111: color_data = 12'b101000000000;
20'b00101101110101010000: color_data = 12'b111000000000;
20'b00101101110101010001: color_data = 12'b111000000000;
20'b00101101110101010010: color_data = 12'b101000000001;
20'b00101101110101010011: color_data = 12'b010100000000;
20'b00101101110101010100: color_data = 12'b001000000000;
20'b00101101110101011111: color_data = 12'b111011101111;
20'b00101101110101100000: color_data = 12'b111011101110;
20'b00101101110101100001: color_data = 12'b111111111110;
20'b00101101110101100010: color_data = 12'b111011101110;
20'b00101101110101100100: color_data = 12'b111011101110;
20'b00101101110101100101: color_data = 12'b111011101110;
20'b00101101110101100110: color_data = 12'b111011101110;
20'b00101101110101100111: color_data = 12'b111011101110;
20'b00101101110101101000: color_data = 12'b111011101110;
20'b00101101110101101111: color_data = 12'b000000010000;
20'b00101101110101110000: color_data = 12'b000000010000;
20'b00101101110101110001: color_data = 12'b000000010000;
20'b00101101110101110010: color_data = 12'b000000010000;
20'b00101101110101110011: color_data = 12'b000000010000;
20'b00101101110101111010: color_data = 12'b111011101110;
20'b00101101110101111011: color_data = 12'b111011101110;
20'b00101101110101111100: color_data = 12'b111011111111;
20'b00101101110101111101: color_data = 12'b111011101110;
20'b00101101110101111110: color_data = 12'b111011101110;
20'b00101101110110000000: color_data = 12'b111011101110;
20'b00101101110110000001: color_data = 12'b111111111111;
20'b00101101110110000010: color_data = 12'b111011101110;
20'b00101101110110000011: color_data = 12'b111011101110;
20'b00101101110110000100: color_data = 12'b111011101110;
20'b00101101110110000110: color_data = 12'b111011101110;
20'b00101101110110000111: color_data = 12'b111111111111;
20'b00101101110110001000: color_data = 12'b111011101110;
20'b00101101110110001001: color_data = 12'b111011101110;
20'b00101101110110001011: color_data = 12'b111011101110;
20'b00101101110110001100: color_data = 12'b111011101110;
20'b00101101110110001101: color_data = 12'b111011101110;
20'b00101101110110001110: color_data = 12'b111011101110;
20'b00101101110110010000: color_data = 12'b111011101110;
20'b00101101110110010001: color_data = 12'b111011101110;
20'b00101101110110010010: color_data = 12'b111111111111;
20'b00101101110110010011: color_data = 12'b111011101110;
20'b00101101110110010100: color_data = 12'b111011101110;
20'b00101110000011110110: color_data = 12'b111111111111;
20'b00101110000011110111: color_data = 12'b111011101110;
20'b00101110000011111000: color_data = 12'b111011101110;
20'b00101110000011111001: color_data = 12'b111011101110;
20'b00101110000011111010: color_data = 12'b111011101110;
20'b00101110000011111100: color_data = 12'b111011101110;
20'b00101110000011111101: color_data = 12'b111011101110;
20'b00101110000011111110: color_data = 12'b111011101110;
20'b00101110000011111111: color_data = 12'b111011101110;
20'b00101110000100000001: color_data = 12'b111011101110;
20'b00101110000100000010: color_data = 12'b111111111111;
20'b00101110000100000011: color_data = 12'b111011101110;
20'b00101110000100000100: color_data = 12'b111011101110;
20'b00101110000100000101: color_data = 12'b111111111111;
20'b00101110000100000111: color_data = 12'b111011101110;
20'b00101110000100001000: color_data = 12'b111011101110;
20'b00101110000100001001: color_data = 12'b111011101110;
20'b00101110000100001010: color_data = 12'b111011101110;
20'b00101110000100001011: color_data = 12'b111011101110;
20'b00101110000100100011: color_data = 12'b111011101110;
20'b00101110000100100100: color_data = 12'b111011101110;
20'b00101110000100100101: color_data = 12'b111011101110;
20'b00101110000100100110: color_data = 12'b111011101110;
20'b00101110000101000111: color_data = 12'b001000000000;
20'b00101110000101001000: color_data = 12'b010100000000;
20'b00101110000101001001: color_data = 12'b101000000000;
20'b00101110000101001010: color_data = 12'b110100000000;
20'b00101110000101001011: color_data = 12'b111000000000;
20'b00101110000101001100: color_data = 12'b111100000000;
20'b00101110000101001101: color_data = 12'b111000000000;
20'b00101110000101001110: color_data = 12'b100100000000;
20'b00101110000101001111: color_data = 12'b101000000000;
20'b00101110000101010000: color_data = 12'b110100000000;
20'b00101110000101010001: color_data = 12'b110100000000;
20'b00101110000101010010: color_data = 12'b101000000001;
20'b00101110000101010011: color_data = 12'b010100000000;
20'b00101110000101010100: color_data = 12'b001000000000;
20'b00101110000101011111: color_data = 12'b111011101110;
20'b00101110000101100000: color_data = 12'b111011111110;
20'b00101110000101100001: color_data = 12'b111011101110;
20'b00101110000101100010: color_data = 12'b111011101110;
20'b00101110000101100100: color_data = 12'b111011101111;
20'b00101110000101100101: color_data = 12'b110111101110;
20'b00101110000101100110: color_data = 12'b111011101110;
20'b00101110000101100111: color_data = 12'b111011111110;
20'b00101110000101101000: color_data = 12'b111011101110;
20'b00101110000101111010: color_data = 12'b111111101110;
20'b00101110000101111011: color_data = 12'b111111101110;
20'b00101110000101111100: color_data = 12'b111111101110;
20'b00101110000101111101: color_data = 12'b111011101110;
20'b00101110000101111110: color_data = 12'b111011101110;
20'b00101110000110000000: color_data = 12'b111011101110;
20'b00101110000110000001: color_data = 12'b111011101110;
20'b00101110000110000010: color_data = 12'b111011101110;
20'b00101110000110000011: color_data = 12'b111111111111;
20'b00101110000110000100: color_data = 12'b111011101110;
20'b00101110000110000110: color_data = 12'b111011101110;
20'b00101110000110000111: color_data = 12'b111011101110;
20'b00101110000110001000: color_data = 12'b111011101110;
20'b00101110000110001001: color_data = 12'b111011101110;
20'b00101110000110001011: color_data = 12'b111011101110;
20'b00101110000110001100: color_data = 12'b111011101110;
20'b00101110000110001101: color_data = 12'b111011101110;
20'b00101110000110001110: color_data = 12'b111011101110;
20'b00101110000110010000: color_data = 12'b111011101110;
20'b00101110000110010001: color_data = 12'b111011101110;
20'b00101110000110010010: color_data = 12'b111111111111;
20'b00101110000110010011: color_data = 12'b111011101110;
20'b00101110000110010100: color_data = 12'b111011101110;
20'b00101110010011110110: color_data = 12'b111011101110;
20'b00101110010011110111: color_data = 12'b111111111111;
20'b00101110010011111000: color_data = 12'b111011101110;
20'b00101110010011111001: color_data = 12'b111011101110;
20'b00101110010011111010: color_data = 12'b111011101110;
20'b00101110010011111100: color_data = 12'b111111111111;
20'b00101110010011111101: color_data = 12'b111111111111;
20'b00101110010011111110: color_data = 12'b111011101110;
20'b00101110010011111111: color_data = 12'b111011101110;
20'b00101110010100000001: color_data = 12'b111011101110;
20'b00101110010100000010: color_data = 12'b111011101110;
20'b00101110010100000011: color_data = 12'b111011101110;
20'b00101110010100000100: color_data = 12'b111011101110;
20'b00101110010100000101: color_data = 12'b111011101110;
20'b00101110010100000111: color_data = 12'b111011101110;
20'b00101110010100001000: color_data = 12'b111011101110;
20'b00101110010100001001: color_data = 12'b111111111111;
20'b00101110010100001010: color_data = 12'b111011101110;
20'b00101110010100001011: color_data = 12'b111011101110;
20'b00101110010100100011: color_data = 12'b111011101110;
20'b00101110010100100100: color_data = 12'b111011101110;
20'b00101110010100100101: color_data = 12'b111111111111;
20'b00101110010100100110: color_data = 12'b111011101110;
20'b00101110010101000111: color_data = 12'b000100000000;
20'b00101110010101001000: color_data = 12'b010000000000;
20'b00101110010101001001: color_data = 12'b100100000000;
20'b00101110010101001010: color_data = 12'b110000000000;
20'b00101110010101001011: color_data = 12'b110100000000;
20'b00101110010101001100: color_data = 12'b111000000000;
20'b00101110010101001101: color_data = 12'b110000000000;
20'b00101110010101001110: color_data = 12'b100000000000;
20'b00101110010101001111: color_data = 12'b100100000000;
20'b00101110010101010000: color_data = 12'b110000000000;
20'b00101110010101010001: color_data = 12'b110000000000;
20'b00101110010101010010: color_data = 12'b100100000000;
20'b00101110010101010011: color_data = 12'b010000000000;
20'b00101110010101010100: color_data = 12'b000100000000;
20'b00101110010101011111: color_data = 12'b111011101110;
20'b00101110010101100000: color_data = 12'b111011101110;
20'b00101110010101100001: color_data = 12'b111011101110;
20'b00101110010101100010: color_data = 12'b111011111111;
20'b00101110010101100100: color_data = 12'b111011101110;
20'b00101110010101100101: color_data = 12'b111011111111;
20'b00101110010101100110: color_data = 12'b111011101110;
20'b00101110010101100111: color_data = 12'b111011101110;
20'b00101110010101101000: color_data = 12'b111011101110;
20'b00101110010101101100: color_data = 12'b000100000000;
20'b00101110010101111010: color_data = 12'b111111101110;
20'b00101110010101111011: color_data = 12'b111011101110;
20'b00101110010101111100: color_data = 12'b111111101110;
20'b00101110010101111101: color_data = 12'b111011101110;
20'b00101110010101111110: color_data = 12'b111011101111;
20'b00101110010110000000: color_data = 12'b111011111111;
20'b00101110010110000001: color_data = 12'b111011101110;
20'b00101110010110000010: color_data = 12'b111011101110;
20'b00101110010110000011: color_data = 12'b111011101110;
20'b00101110010110000100: color_data = 12'b111111111111;
20'b00101110010110000110: color_data = 12'b111011101110;
20'b00101110010110000111: color_data = 12'b111011101110;
20'b00101110010110001000: color_data = 12'b111011101110;
20'b00101110010110001001: color_data = 12'b111011101110;
20'b00101110010110001011: color_data = 12'b111011101110;
20'b00101110010110001100: color_data = 12'b111011101110;
20'b00101110010110001101: color_data = 12'b111011101110;
20'b00101110010110001110: color_data = 12'b111011101110;
20'b00101110010110010000: color_data = 12'b111111111111;
20'b00101110010110010001: color_data = 12'b111111111111;
20'b00101110010110010010: color_data = 12'b111011101110;
20'b00101110010110010011: color_data = 12'b111011101110;
20'b00101110010110010100: color_data = 12'b111011101110;
20'b00101110100011110110: color_data = 12'b111111111111;
20'b00101110100011110111: color_data = 12'b111011101110;
20'b00101110100011111000: color_data = 12'b111111111111;
20'b00101110100011111001: color_data = 12'b111011101110;
20'b00101110100011111010: color_data = 12'b111011101110;
20'b00101110100011111100: color_data = 12'b111011101110;
20'b00101110100011111101: color_data = 12'b111011101110;
20'b00101110100011111110: color_data = 12'b111011101110;
20'b00101110100011111111: color_data = 12'b111011101110;
20'b00101110100100000001: color_data = 12'b111111111111;
20'b00101110100100000010: color_data = 12'b111011101110;
20'b00101110100100000011: color_data = 12'b111011101110;
20'b00101110100100000100: color_data = 12'b111011101110;
20'b00101110100100000101: color_data = 12'b111011101110;
20'b00101110100100000111: color_data = 12'b111011101110;
20'b00101110100100001000: color_data = 12'b111011101110;
20'b00101110100100001001: color_data = 12'b111011101110;
20'b00101110100100001010: color_data = 12'b111011101110;
20'b00101110100100001011: color_data = 12'b111111111111;
20'b00101110100100100011: color_data = 12'b111011101110;
20'b00101110100100100100: color_data = 12'b111011101110;
20'b00101110100100100101: color_data = 12'b111011101110;
20'b00101110100100100110: color_data = 12'b111011101110;
20'b00101110100101001000: color_data = 12'b001100000000;
20'b00101110100101001001: color_data = 12'b011100000001;
20'b00101110100101001010: color_data = 12'b100100000001;
20'b00101110100101001011: color_data = 12'b101000000000;
20'b00101110100101001100: color_data = 12'b101000000000;
20'b00101110100101001101: color_data = 12'b100100000000;
20'b00101110100101001110: color_data = 12'b011000000000;
20'b00101110100101001111: color_data = 12'b011100000001;
20'b00101110100101010000: color_data = 12'b100100010001;
20'b00101110100101010001: color_data = 12'b100100000000;
20'b00101110100101010010: color_data = 12'b011100010001;
20'b00101110100101010011: color_data = 12'b001100000000;
20'b00101110100101010100: color_data = 12'b000100000000;
20'b00101110100101011111: color_data = 12'b111011101110;
20'b00101110100101100000: color_data = 12'b111011101110;
20'b00101110100101100001: color_data = 12'b111011111110;
20'b00101110100101100010: color_data = 12'b111011101110;
20'b00101110100101100100: color_data = 12'b111011101111;
20'b00101110100101100101: color_data = 12'b111011101110;
20'b00101110100101100110: color_data = 12'b111111111110;
20'b00101110100101100111: color_data = 12'b111111101110;
20'b00101110100101101000: color_data = 12'b111011101110;
20'b00101110100101111010: color_data = 12'b111011101110;
20'b00101110100101111011: color_data = 12'b111111101110;
20'b00101110100101111100: color_data = 12'b111111111111;
20'b00101110100101111101: color_data = 12'b111011101110;
20'b00101110100101111110: color_data = 12'b111111111110;
20'b00101110100110000000: color_data = 12'b111011101110;
20'b00101110100110000001: color_data = 12'b111011101110;
20'b00101110100110000010: color_data = 12'b111011101110;
20'b00101110100110000011: color_data = 12'b111011101110;
20'b00101110100110000100: color_data = 12'b111011101110;
20'b00101110100110000110: color_data = 12'b111011101110;
20'b00101110100110000111: color_data = 12'b111111111111;
20'b00101110100110001000: color_data = 12'b111011101110;
20'b00101110100110001001: color_data = 12'b111011101110;
20'b00101110100110001011: color_data = 12'b111011101110;
20'b00101110100110001100: color_data = 12'b111011101110;
20'b00101110100110001101: color_data = 12'b111011101110;
20'b00101110100110001110: color_data = 12'b111011101110;
20'b00101110100110010000: color_data = 12'b111011101110;
20'b00101110100110010001: color_data = 12'b111011101110;
20'b00101110100110010010: color_data = 12'b111111111111;
20'b00101110100110010011: color_data = 12'b111011101110;
20'b00101110100110010100: color_data = 12'b111011101110;
20'b00101110110101001000: color_data = 12'b000100000000;
20'b00101110110101001001: color_data = 12'b001100000000;
20'b00101110110101001010: color_data = 12'b010100000000;
20'b00101110110101001011: color_data = 12'b010100000000;
20'b00101110110101001100: color_data = 12'b010100000000;
20'b00101110110101001101: color_data = 12'b010100000000;
20'b00101110110101001110: color_data = 12'b001100000000;
20'b00101110110101001111: color_data = 12'b001100000000;
20'b00101110110101010000: color_data = 12'b010000000000;
20'b00101110110101010001: color_data = 12'b010000000000;
20'b00101110110101010010: color_data = 12'b001100000000;
20'b00101110110101010011: color_data = 12'b001000000000;
20'b00101111000100000111: color_data = 12'b111011101110;
20'b00101111000100001000: color_data = 12'b111011101110;
20'b00101111000100001001: color_data = 12'b111011101110;
20'b00101111000100001010: color_data = 12'b111011101110;
20'b00101111000100001011: color_data = 12'b111011101110;
20'b00101111000100001101: color_data = 12'b111011101110;
20'b00101111000100001110: color_data = 12'b111011101110;
20'b00101111000100001111: color_data = 12'b111111111111;
20'b00101111000100010000: color_data = 12'b111011101110;
20'b00101111000100011101: color_data = 12'b111111111111;
20'b00101111000100011110: color_data = 12'b111011101110;
20'b00101111000100011111: color_data = 12'b111111111111;
20'b00101111000100100000: color_data = 12'b111011101110;
20'b00101111000100100001: color_data = 12'b111011101110;
20'b00101111000100100011: color_data = 12'b111011101110;
20'b00101111000100100100: color_data = 12'b111011101110;
20'b00101111000100100101: color_data = 12'b111011101110;
20'b00101111000100100110: color_data = 12'b111011101110;
20'b00101111000100110011: color_data = 12'b111011101110;
20'b00101111000100110100: color_data = 12'b111111111111;
20'b00101111000100110101: color_data = 12'b111011101110;
20'b00101111000100110110: color_data = 12'b111011101110;
20'b00101111000100110111: color_data = 12'b111011101110;
20'b00101111000101000011: color_data = 12'b111011101110;
20'b00101111000101000100: color_data = 12'b111011111111;
20'b00101111000101000101: color_data = 12'b111011101110;
20'b00101111000101000110: color_data = 12'b111011101110;
20'b00101111000101000111: color_data = 12'b111111101110;
20'b00101111000101001010: color_data = 12'b000100000000;
20'b00101111000101001011: color_data = 12'b000100000000;
20'b00101111000101001100: color_data = 12'b000100000000;
20'b00101111000101001101: color_data = 12'b000100000000;
20'b00101111000101001111: color_data = 12'b000100000000;
20'b00101111000101010000: color_data = 12'b000100000000;
20'b00101111000101010001: color_data = 12'b000100000000;
20'b00101111000101010010: color_data = 12'b000100000000;
20'b00101111000101010011: color_data = 12'b000100000000;
20'b00101111000101011001: color_data = 12'b111011101110;
20'b00101111000101011010: color_data = 12'b111011101110;
20'b00101111000101011011: color_data = 12'b111011101110;
20'b00101111000101011100: color_data = 12'b111111101110;
20'b00101111000101011101: color_data = 12'b111111101110;
20'b00101111000101011111: color_data = 12'b111011101110;
20'b00101111000101100000: color_data = 12'b111011101110;
20'b00101111000101100001: color_data = 12'b111011101110;
20'b00101111000101100010: color_data = 12'b111011101110;
20'b00101111000101100100: color_data = 12'b111011101111;
20'b00101111000101100101: color_data = 12'b111011101110;
20'b00101111000101100110: color_data = 12'b111111111111;
20'b00101111000101100111: color_data = 12'b111011101110;
20'b00101111000101101000: color_data = 12'b111111111110;
20'b00101111000101110101: color_data = 12'b111011111111;
20'b00101111000101110110: color_data = 12'b111011101110;
20'b00101111000101110111: color_data = 12'b111011111110;
20'b00101111000101111000: color_data = 12'b111011111111;
20'b00101111000101111001: color_data = 12'b111011101110;
20'b00101111010100000111: color_data = 12'b111111111111;
20'b00101111010100001000: color_data = 12'b111011101110;
20'b00101111010100001001: color_data = 12'b111011101110;
20'b00101111010100001010: color_data = 12'b111011101110;
20'b00101111010100001011: color_data = 12'b111011101110;
20'b00101111010100001101: color_data = 12'b111111111111;
20'b00101111010100001110: color_data = 12'b111011101110;
20'b00101111010100001111: color_data = 12'b111011101110;
20'b00101111010100010000: color_data = 12'b111011101110;
20'b00101111010100011101: color_data = 12'b111011101110;
20'b00101111010100011110: color_data = 12'b111011101110;
20'b00101111010100011111: color_data = 12'b111011101110;
20'b00101111010100100000: color_data = 12'b111111111111;
20'b00101111010100100001: color_data = 12'b111011101110;
20'b00101111010100100011: color_data = 12'b111011101110;
20'b00101111010100100100: color_data = 12'b111011101110;
20'b00101111010100100101: color_data = 12'b111011101110;
20'b00101111010100100110: color_data = 12'b111011101110;
20'b00101111010100110011: color_data = 12'b111111111111;
20'b00101111010100110100: color_data = 12'b111011101110;
20'b00101111010100110101: color_data = 12'b111011101110;
20'b00101111010100110110: color_data = 12'b111011101110;
20'b00101111010100110111: color_data = 12'b111011101110;
20'b00101111010101000011: color_data = 12'b111011101111;
20'b00101111010101000100: color_data = 12'b111011101110;
20'b00101111010101000101: color_data = 12'b111011101110;
20'b00101111010101000110: color_data = 12'b111011101110;
20'b00101111010101000111: color_data = 12'b111111101110;
20'b00101111010101011001: color_data = 12'b111011101111;
20'b00101111010101011010: color_data = 12'b111011101110;
20'b00101111010101011011: color_data = 12'b111011101111;
20'b00101111010101011100: color_data = 12'b111011101110;
20'b00101111010101011101: color_data = 12'b111011101110;
20'b00101111010101011111: color_data = 12'b111111101110;
20'b00101111010101100000: color_data = 12'b111011101110;
20'b00101111010101100001: color_data = 12'b111111111110;
20'b00101111010101100010: color_data = 12'b111011101110;
20'b00101111010101100100: color_data = 12'b111011101110;
20'b00101111010101100101: color_data = 12'b111011111111;
20'b00101111010101100110: color_data = 12'b111011101110;
20'b00101111010101100111: color_data = 12'b111011101110;
20'b00101111010101101000: color_data = 12'b111011101110;
20'b00101111010101110101: color_data = 12'b111011101110;
20'b00101111010101110110: color_data = 12'b111011101110;
20'b00101111010101110111: color_data = 12'b111011101110;
20'b00101111010101111000: color_data = 12'b111011101110;
20'b00101111010101111001: color_data = 12'b111011101110;
20'b00101111100100000111: color_data = 12'b111011101110;
20'b00101111100100001000: color_data = 12'b111011101110;
20'b00101111100100001001: color_data = 12'b111011101110;
20'b00101111100100001010: color_data = 12'b111011101110;
20'b00101111100100001011: color_data = 12'b111011101110;
20'b00101111100100001101: color_data = 12'b111011101110;
20'b00101111100100001110: color_data = 12'b111011101110;
20'b00101111100100001111: color_data = 12'b111011101110;
20'b00101111100100010000: color_data = 12'b111011101110;
20'b00101111100100011101: color_data = 12'b111011101110;
20'b00101111100100011110: color_data = 12'b111011101110;
20'b00101111100100011111: color_data = 12'b111011101110;
20'b00101111100100100000: color_data = 12'b111011101110;
20'b00101111100100100001: color_data = 12'b111011101110;
20'b00101111100100100011: color_data = 12'b111111111111;
20'b00101111100100100100: color_data = 12'b111011101110;
20'b00101111100100100101: color_data = 12'b111011101110;
20'b00101111100100100110: color_data = 12'b111011101110;
20'b00101111100100110011: color_data = 12'b111011101110;
20'b00101111100100110100: color_data = 12'b111011101110;
20'b00101111100100110101: color_data = 12'b111011101110;
20'b00101111100100110110: color_data = 12'b111011101110;
20'b00101111100100110111: color_data = 12'b111011101110;
20'b00101111100101000011: color_data = 12'b111011101111;
20'b00101111100101000100: color_data = 12'b111011101110;
20'b00101111100101000101: color_data = 12'b111011111110;
20'b00101111100101000110: color_data = 12'b111011111110;
20'b00101111100101000111: color_data = 12'b111011101110;
20'b00101111100101011001: color_data = 12'b111011101110;
20'b00101111100101011010: color_data = 12'b111111101111;
20'b00101111100101011011: color_data = 12'b111111101111;
20'b00101111100101011100: color_data = 12'b111011101110;
20'b00101111100101011101: color_data = 12'b111111111111;
20'b00101111100101011111: color_data = 12'b111011101110;
20'b00101111100101100000: color_data = 12'b111011101110;
20'b00101111100101100001: color_data = 12'b111011101110;
20'b00101111100101100010: color_data = 12'b111011101110;
20'b00101111100101100100: color_data = 12'b111011101111;
20'b00101111100101100101: color_data = 12'b111011101110;
20'b00101111100101100110: color_data = 12'b111011101110;
20'b00101111100101100111: color_data = 12'b111011111110;
20'b00101111100101101000: color_data = 12'b111011101110;
20'b00101111100101110101: color_data = 12'b111011101110;
20'b00101111100101110110: color_data = 12'b111011101110;
20'b00101111100101110111: color_data = 12'b111011101110;
20'b00101111100101111000: color_data = 12'b111011101110;
20'b00101111100101111001: color_data = 12'b111011101110;
20'b00101111110100000111: color_data = 12'b111011101110;
20'b00101111110100001000: color_data = 12'b111111111111;
20'b00101111110100001001: color_data = 12'b111011101110;
20'b00101111110100001010: color_data = 12'b111011101110;
20'b00101111110100001011: color_data = 12'b111111111111;
20'b00101111110100001101: color_data = 12'b111011101110;
20'b00101111110100001110: color_data = 12'b111111111111;
20'b00101111110100001111: color_data = 12'b111011101110;
20'b00101111110100010000: color_data = 12'b111011101110;
20'b00101111110100011101: color_data = 12'b111011101110;
20'b00101111110100011110: color_data = 12'b111011101110;
20'b00101111110100011111: color_data = 12'b111011101110;
20'b00101111110100100000: color_data = 12'b111011101110;
20'b00101111110100100001: color_data = 12'b111011101110;
20'b00101111110100100011: color_data = 12'b111011101110;
20'b00101111110100100100: color_data = 12'b111011101110;
20'b00101111110100100101: color_data = 12'b111011101110;
20'b00101111110100100110: color_data = 12'b111011101110;
20'b00101111110100110011: color_data = 12'b111011101110;
20'b00101111110100110100: color_data = 12'b111011101110;
20'b00101111110100110101: color_data = 12'b111011101110;
20'b00101111110100110110: color_data = 12'b111011101110;
20'b00101111110100110111: color_data = 12'b111011101110;
20'b00101111110101000011: color_data = 12'b111011101110;
20'b00101111110101000100: color_data = 12'b111011101110;
20'b00101111110101000101: color_data = 12'b111011101110;
20'b00101111110101000110: color_data = 12'b111011101110;
20'b00101111110101000111: color_data = 12'b111011101110;
20'b00101111110101011001: color_data = 12'b111111101111;
20'b00101111110101011010: color_data = 12'b111011101110;
20'b00101111110101011011: color_data = 12'b111011101110;
20'b00101111110101011100: color_data = 12'b111011101110;
20'b00101111110101011101: color_data = 12'b111011101110;
20'b00101111110101011111: color_data = 12'b111011101110;
20'b00101111110101100000: color_data = 12'b111011101110;
20'b00101111110101100001: color_data = 12'b111011101110;
20'b00101111110101100010: color_data = 12'b111011101110;
20'b00101111110101100100: color_data = 12'b111011101110;
20'b00101111110101100101: color_data = 12'b111011101110;
20'b00101111110101100110: color_data = 12'b111011111110;
20'b00101111110101100111: color_data = 12'b111011101110;
20'b00101111110101101000: color_data = 12'b111011101110;
20'b00101111110101110101: color_data = 12'b111011101110;
20'b00101111110101110110: color_data = 12'b111011101110;
20'b00101111110101110111: color_data = 12'b111111111110;
20'b00101111110101111000: color_data = 12'b111011111110;
20'b00101111110101111001: color_data = 12'b111011101110;
20'b00110000000100000111: color_data = 12'b111011101110;
20'b00110000000100001000: color_data = 12'b111011101110;
20'b00110000000100001001: color_data = 12'b111011101110;
20'b00110000000100001010: color_data = 12'b111011101110;
20'b00110000000100001011: color_data = 12'b111011101110;
20'b00110000000100001101: color_data = 12'b111011101110;
20'b00110000000100001110: color_data = 12'b111011101110;
20'b00110000000100001111: color_data = 12'b111011101110;
20'b00110000000100010000: color_data = 12'b111011101110;
20'b00110000010011101011: color_data = 12'b111011101110;
20'b00110000010011101100: color_data = 12'b111011101110;
20'b00110000010011101101: color_data = 12'b111011101110;
20'b00110000010011101110: color_data = 12'b111011101110;
20'b00110000010011101111: color_data = 12'b111011101110;
20'b00110000010011110001: color_data = 12'b111011101110;
20'b00110000010011110010: color_data = 12'b111011101110;
20'b00110000010011110011: color_data = 12'b111011101110;
20'b00110000010011110100: color_data = 12'b111011101110;
20'b00110000010011110101: color_data = 12'b111111111111;
20'b00110000010100010111: color_data = 12'b111011101110;
20'b00110000010100011000: color_data = 12'b111111111111;
20'b00110000010100011001: color_data = 12'b111111111111;
20'b00110000010100011010: color_data = 12'b111011101110;
20'b00110000010100011011: color_data = 12'b111011101110;
20'b00110000010100011101: color_data = 12'b111011101110;
20'b00110000010100011110: color_data = 12'b111011101110;
20'b00110000010100011111: color_data = 12'b111011101110;
20'b00110000010100100000: color_data = 12'b111011101110;
20'b00110000010100100001: color_data = 12'b111111111111;
20'b00110000010100110011: color_data = 12'b111011101110;
20'b00110000010100110100: color_data = 12'b111011101110;
20'b00110000010100110101: color_data = 12'b111011101110;
20'b00110000010100110110: color_data = 12'b111011101110;
20'b00110000010100110111: color_data = 12'b111011101110;
20'b00110000010100111001: color_data = 12'b111011101110;
20'b00110000010100111010: color_data = 12'b111011101110;
20'b00110000010100111011: color_data = 12'b111011101110;
20'b00110000010100111100: color_data = 12'b111011101110;
20'b00110000010101000011: color_data = 12'b111011101110;
20'b00110000010101000100: color_data = 12'b111011101110;
20'b00110000010101000101: color_data = 12'b111011101110;
20'b00110000010101000110: color_data = 12'b111011101110;
20'b00110000010101000111: color_data = 12'b111011101110;
20'b00110000010101001001: color_data = 12'b111011101110;
20'b00110000010101001010: color_data = 12'b111111111111;
20'b00110000010101001011: color_data = 12'b111011101110;
20'b00110000010101001100: color_data = 12'b111011101110;
20'b00110000010101001101: color_data = 12'b111011101110;
20'b00110000010101001111: color_data = 12'b111011101110;
20'b00110000010101010000: color_data = 12'b111011101110;
20'b00110000010101010001: color_data = 12'b111011101110;
20'b00110000010101010010: color_data = 12'b111011101110;
20'b00110000010101010100: color_data = 12'b111011101110;
20'b00110000010101010101: color_data = 12'b111011101110;
20'b00110000010101010110: color_data = 12'b111011101110;
20'b00110000010101010111: color_data = 12'b111011101110;
20'b00110000010101011001: color_data = 12'b111111111111;
20'b00110000010101011010: color_data = 12'b111011101110;
20'b00110000010101011011: color_data = 12'b111011101110;
20'b00110000010101011100: color_data = 12'b111011101110;
20'b00110000010101011101: color_data = 12'b111011101110;
20'b00110000010101011111: color_data = 12'b111011101110;
20'b00110000010101100000: color_data = 12'b111011101110;
20'b00110000010101100001: color_data = 12'b111011101110;
20'b00110000010101100010: color_data = 12'b111011101110;
20'b00110000010101100100: color_data = 12'b111011101110;
20'b00110000010101100101: color_data = 12'b111011101110;
20'b00110000010101100110: color_data = 12'b111111111111;
20'b00110000010101100111: color_data = 12'b111111111111;
20'b00110000010101101000: color_data = 12'b111011101110;
20'b00110000010101110101: color_data = 12'b111011101110;
20'b00110000010101110110: color_data = 12'b111011101110;
20'b00110000010101110111: color_data = 12'b111011101110;
20'b00110000010101111000: color_data = 12'b111011101110;
20'b00110000010101111001: color_data = 12'b111011101110;
20'b00110000100011101011: color_data = 12'b111011101110;
20'b00110000100011101100: color_data = 12'b111011101110;
20'b00110000100011101101: color_data = 12'b111011101110;
20'b00110000100011101110: color_data = 12'b111011101110;
20'b00110000100011101111: color_data = 12'b111011101110;
20'b00110000100011110001: color_data = 12'b111011101110;
20'b00110000100011110010: color_data = 12'b111011101110;
20'b00110000100011110011: color_data = 12'b111111111111;
20'b00110000100011110100: color_data = 12'b111111111111;
20'b00110000100011110101: color_data = 12'b111011101110;
20'b00110000100100010111: color_data = 12'b111011101110;
20'b00110000100100011000: color_data = 12'b111011101110;
20'b00110000100100011001: color_data = 12'b111011101110;
20'b00110000100100011010: color_data = 12'b111011101110;
20'b00110000100100011011: color_data = 12'b111011101110;
20'b00110000100100011101: color_data = 12'b111011101110;
20'b00110000100100011110: color_data = 12'b111111111111;
20'b00110000100100011111: color_data = 12'b111011101110;
20'b00110000100100100000: color_data = 12'b111011101110;
20'b00110000100100100001: color_data = 12'b111011101110;
20'b00110000100100110011: color_data = 12'b111011101110;
20'b00110000100100110100: color_data = 12'b111011101110;
20'b00110000100100110101: color_data = 12'b111011101110;
20'b00110000100100110110: color_data = 12'b111011101110;
20'b00110000100100110111: color_data = 12'b111011101110;
20'b00110000100100111001: color_data = 12'b111011101110;
20'b00110000100100111010: color_data = 12'b111011101110;
20'b00110000100100111011: color_data = 12'b111011101110;
20'b00110000100100111100: color_data = 12'b111111111111;
20'b00110000100101000011: color_data = 12'b111011101110;
20'b00110000100101000100: color_data = 12'b111011101110;
20'b00110000100101000101: color_data = 12'b111011101110;
20'b00110000100101000110: color_data = 12'b111011101110;
20'b00110000100101000111: color_data = 12'b111011101110;
20'b00110000100101001001: color_data = 12'b111011101110;
20'b00110000100101001010: color_data = 12'b111011101110;
20'b00110000100101001011: color_data = 12'b111011101110;
20'b00110000100101001100: color_data = 12'b111011101110;
20'b00110000100101001101: color_data = 12'b111011101110;
20'b00110000100101001111: color_data = 12'b111011101110;
20'b00110000100101010000: color_data = 12'b111011101110;
20'b00110000100101010001: color_data = 12'b111011101110;
20'b00110000100101010010: color_data = 12'b111011101110;
20'b00110000100101010100: color_data = 12'b111011101110;
20'b00110000100101010101: color_data = 12'b111011101110;
20'b00110000100101010110: color_data = 12'b111111111111;
20'b00110000100101010111: color_data = 12'b111011101110;
20'b00110000100101011001: color_data = 12'b111011101110;
20'b00110000100101011010: color_data = 12'b111011101110;
20'b00110000100101011011: color_data = 12'b111011101110;
20'b00110000100101011100: color_data = 12'b111011101110;
20'b00110000100101011101: color_data = 12'b111011101110;
20'b00110000100101011111: color_data = 12'b111011101110;
20'b00110000100101100000: color_data = 12'b111011101110;
20'b00110000100101100001: color_data = 12'b111111111111;
20'b00110000100101100010: color_data = 12'b111011101110;
20'b00110000100101100100: color_data = 12'b111011101110;
20'b00110000100101100101: color_data = 12'b111011101110;
20'b00110000100101100110: color_data = 12'b111011101110;
20'b00110000100101100111: color_data = 12'b111011101110;
20'b00110000100101101000: color_data = 12'b111011101110;
20'b00110000100101110101: color_data = 12'b111011101110;
20'b00110000100101110110: color_data = 12'b111011101110;
20'b00110000100101110111: color_data = 12'b111011101110;
20'b00110000100101111000: color_data = 12'b111011101110;
20'b00110000100101111001: color_data = 12'b111011101110;
20'b00110000110011101011: color_data = 12'b111111111111;
20'b00110000110011101100: color_data = 12'b111011101110;
20'b00110000110011101101: color_data = 12'b111011101110;
20'b00110000110011101110: color_data = 12'b111011101110;
20'b00110000110011101111: color_data = 12'b111011101110;
20'b00110000110011110001: color_data = 12'b111011101110;
20'b00110000110011110010: color_data = 12'b111111111111;
20'b00110000110011110011: color_data = 12'b111011101110;
20'b00110000110011110100: color_data = 12'b111011101110;
20'b00110000110011110101: color_data = 12'b111011101110;
20'b00110000110100010111: color_data = 12'b111011101110;
20'b00110000110100011000: color_data = 12'b111011101110;
20'b00110000110100011001: color_data = 12'b111111111111;
20'b00110000110100011010: color_data = 12'b111111111111;
20'b00110000110100011011: color_data = 12'b111011101110;
20'b00110000110100011101: color_data = 12'b111011101110;
20'b00110000110100011110: color_data = 12'b111011101110;
20'b00110000110100011111: color_data = 12'b111011101110;
20'b00110000110100100000: color_data = 12'b111111111111;
20'b00110000110100100001: color_data = 12'b111011101110;
20'b00110000110100110011: color_data = 12'b111111111111;
20'b00110000110100110100: color_data = 12'b111011101110;
20'b00110000110100110101: color_data = 12'b111011101110;
20'b00110000110100110110: color_data = 12'b111011101110;
20'b00110000110100110111: color_data = 12'b111011101110;
20'b00110000110100111001: color_data = 12'b111011101110;
20'b00110000110100111010: color_data = 12'b111011101110;
20'b00110000110100111011: color_data = 12'b111011101110;
20'b00110000110100111100: color_data = 12'b111011101110;
20'b00110000110101000011: color_data = 12'b111111111111;
20'b00110000110101000100: color_data = 12'b111011101110;
20'b00110000110101000101: color_data = 12'b111011101110;
20'b00110000110101000110: color_data = 12'b111011101110;
20'b00110000110101000111: color_data = 12'b111011101110;
20'b00110000110101001001: color_data = 12'b111011101110;
20'b00110000110101001010: color_data = 12'b111011101110;
20'b00110000110101001011: color_data = 12'b111011101110;
20'b00110000110101001100: color_data = 12'b111011101110;
20'b00110000110101001101: color_data = 12'b111011101110;
20'b00110000110101001111: color_data = 12'b111011101110;
20'b00110000110101010000: color_data = 12'b111011101110;
20'b00110000110101010001: color_data = 12'b111011101110;
20'b00110000110101010010: color_data = 12'b111011101110;
20'b00110000110101010100: color_data = 12'b111011101110;
20'b00110000110101010101: color_data = 12'b111011101110;
20'b00110000110101010110: color_data = 12'b111011101110;
20'b00110000110101010111: color_data = 12'b111011101110;
20'b00110000110101011001: color_data = 12'b111111111111;
20'b00110000110101011010: color_data = 12'b111011101110;
20'b00110000110101011011: color_data = 12'b111011101110;
20'b00110000110101011100: color_data = 12'b111011101110;
20'b00110000110101011101: color_data = 12'b111011101110;
20'b00110000110101011111: color_data = 12'b111011101110;
20'b00110000110101100000: color_data = 12'b111011101110;
20'b00110000110101100001: color_data = 12'b111011101110;
20'b00110000110101100010: color_data = 12'b111011101110;
20'b00110000110101100100: color_data = 12'b111011101110;
20'b00110000110101100101: color_data = 12'b111111111111;
20'b00110000110101100110: color_data = 12'b111111111111;
20'b00110000110101100111: color_data = 12'b111011101110;
20'b00110000110101101000: color_data = 12'b111011101110;
20'b00110000110101110101: color_data = 12'b111011101110;
20'b00110000110101110110: color_data = 12'b111111111111;
20'b00110000110101110111: color_data = 12'b111011101110;
20'b00110000110101111000: color_data = 12'b111011101110;
20'b00110000110101111001: color_data = 12'b111011101110;
20'b00110001000011101011: color_data = 12'b111011101110;
20'b00110001000011101100: color_data = 12'b111011101110;
20'b00110001000011101101: color_data = 12'b111111111111;
20'b00110001000011101110: color_data = 12'b111011101110;
20'b00110001000011101111: color_data = 12'b111011101110;
20'b00110001000011110001: color_data = 12'b111011101110;
20'b00110001000011110010: color_data = 12'b111011101110;
20'b00110001000011110011: color_data = 12'b111011101110;
20'b00110001000011110100: color_data = 12'b111011101110;
20'b00110001000011110101: color_data = 12'b111011101110;
20'b00110001000100010111: color_data = 12'b111011101110;
20'b00110001000100011000: color_data = 12'b111011101110;
20'b00110001000100011001: color_data = 12'b111011101110;
20'b00110001000100011010: color_data = 12'b111011101110;
20'b00110001000100011011: color_data = 12'b111011101110;
20'b00110001000100011101: color_data = 12'b111011101110;
20'b00110001000100011110: color_data = 12'b111011101110;
20'b00110001000100011111: color_data = 12'b111011101110;
20'b00110001000100100000: color_data = 12'b111011101110;
20'b00110001000100100001: color_data = 12'b111111111111;
20'b00110001000100110011: color_data = 12'b111011101110;
20'b00110001000100110100: color_data = 12'b111011101110;
20'b00110001000100110101: color_data = 12'b111111111111;
20'b00110001000100110110: color_data = 12'b111011101110;
20'b00110001000100110111: color_data = 12'b111011101110;
20'b00110001000100111001: color_data = 12'b111011101110;
20'b00110001000100111010: color_data = 12'b111011101110;
20'b00110001000100111011: color_data = 12'b111011101110;
20'b00110001000100111100: color_data = 12'b111011101110;
20'b00110001000101000011: color_data = 12'b111011101110;
20'b00110001000101000100: color_data = 12'b111011101110;
20'b00110001000101000101: color_data = 12'b111111111111;
20'b00110001000101000110: color_data = 12'b111011101110;
20'b00110001000101000111: color_data = 12'b111011101110;
20'b00110001000101001001: color_data = 12'b111011101110;
20'b00110001000101001010: color_data = 12'b111011101110;
20'b00110001000101001011: color_data = 12'b111011101110;
20'b00110001000101001100: color_data = 12'b111011101110;
20'b00110001000101001101: color_data = 12'b111111111111;
20'b00110001000101001111: color_data = 12'b111011101110;
20'b00110001000101010000: color_data = 12'b111011101110;
20'b00110001000101010001: color_data = 12'b111011101110;
20'b00110001000101010010: color_data = 12'b111111111111;
20'b00110001000101010100: color_data = 12'b111011101110;
20'b00110001000101010101: color_data = 12'b111011101110;
20'b00110001000101010110: color_data = 12'b111111111111;
20'b00110001000101010111: color_data = 12'b111011101110;
20'b00110001000101011001: color_data = 12'b111011101110;
20'b00110001000101011010: color_data = 12'b111011101110;
20'b00110001000101011011: color_data = 12'b111011101110;
20'b00110001000101011100: color_data = 12'b111011101110;
20'b00110001000101011101: color_data = 12'b111011101110;
20'b00110001000101011111: color_data = 12'b111111111111;
20'b00110001000101100000: color_data = 12'b111011101110;
20'b00110001000101100001: color_data = 12'b111011101110;
20'b00110001000101100010: color_data = 12'b111011101110;
20'b00110001000101100100: color_data = 12'b111011101110;
20'b00110001000101100101: color_data = 12'b111011101110;
20'b00110001000101100110: color_data = 12'b111011101110;
20'b00110001000101100111: color_data = 12'b111011101110;
20'b00110001000101101000: color_data = 12'b111011101110;
20'b00110001000101110101: color_data = 12'b111011101110;
20'b00110001000101110110: color_data = 12'b111011101110;
20'b00110001000101110111: color_data = 12'b111011101110;
20'b00110001000101111000: color_data = 12'b111011101110;
20'b00110001000101111001: color_data = 12'b111011101110;
20'b00110001100011101011: color_data = 12'b111011101110;
20'b00110001100011101100: color_data = 12'b111011101110;
20'b00110001100011101101: color_data = 12'b111011101110;
20'b00110001100011101110: color_data = 12'b111111111111;
20'b00110001100011101111: color_data = 12'b111011101110;
20'b00110001100011110001: color_data = 12'b111011101110;
20'b00110001100011110010: color_data = 12'b111011101110;
20'b00110001100011110011: color_data = 12'b111011101110;
20'b00110001100011110100: color_data = 12'b111011101110;
20'b00110001100011110101: color_data = 12'b111011101110;
20'b00110001100100010111: color_data = 12'b111011101110;
20'b00110001100100011000: color_data = 12'b111011101110;
20'b00110001100100011001: color_data = 12'b111011101110;
20'b00110001100100011010: color_data = 12'b111011101110;
20'b00110001100100011011: color_data = 12'b111011101110;
20'b00110001100100011101: color_data = 12'b111111111111;
20'b00110001100100011110: color_data = 12'b111011101110;
20'b00110001100100011111: color_data = 12'b111111111111;
20'b00110001100100100000: color_data = 12'b111011101110;
20'b00110001100100100001: color_data = 12'b111011101110;
20'b00110001100100110011: color_data = 12'b111011101110;
20'b00110001100100110100: color_data = 12'b111011101110;
20'b00110001100100110101: color_data = 12'b111011101110;
20'b00110001100100110110: color_data = 12'b111111111111;
20'b00110001100100110111: color_data = 12'b111011101110;
20'b00110001100100111001: color_data = 12'b111011101110;
20'b00110001100100111010: color_data = 12'b111011101110;
20'b00110001100100111011: color_data = 12'b111011101110;
20'b00110001100100111100: color_data = 12'b111111111111;
20'b00110001100101000011: color_data = 12'b111011101110;
20'b00110001100101000100: color_data = 12'b111011101110;
20'b00110001100101000101: color_data = 12'b111011101110;
20'b00110001100101000110: color_data = 12'b111111111111;
20'b00110001100101000111: color_data = 12'b111011101110;
20'b00110001100101001001: color_data = 12'b111011101110;
20'b00110001100101001010: color_data = 12'b111011101110;
20'b00110001100101001011: color_data = 12'b111111111111;
20'b00110001100101001100: color_data = 12'b111011101110;
20'b00110001100101001101: color_data = 12'b111011101110;
20'b00110001100101010100: color_data = 12'b111111111111;
20'b00110001100101010101: color_data = 12'b111011101110;
20'b00110001100101010110: color_data = 12'b111011101110;
20'b00110001100101010111: color_data = 12'b111011101110;
20'b00110001100101011111: color_data = 12'b111011101110;
20'b00110001100101100000: color_data = 12'b111111111111;
20'b00110001100101100001: color_data = 12'b111011101110;
20'b00110001100101100010: color_data = 12'b111111111111;
20'b00110001100101100100: color_data = 12'b111011101110;
20'b00110001100101100101: color_data = 12'b111011101110;
20'b00110001100101100110: color_data = 12'b111011101110;
20'b00110001100101100111: color_data = 12'b111011101110;
20'b00110001100101101000: color_data = 12'b111011101110;
20'b00110001100101101111: color_data = 12'b111011101110;
20'b00110001100101110000: color_data = 12'b111111111111;
20'b00110001100101110001: color_data = 12'b111011101110;
20'b00110001100101110010: color_data = 12'b111011101110;
20'b00110001100101110011: color_data = 12'b111011101110;
20'b00110001100101110101: color_data = 12'b111011101110;
20'b00110001100101110110: color_data = 12'b111011101110;
20'b00110001100101110111: color_data = 12'b111011101110;
20'b00110001100101111000: color_data = 12'b111111111111;
20'b00110001100101111001: color_data = 12'b111011101110;
20'b00110001100101111011: color_data = 12'b111011101110;
20'b00110001100101111100: color_data = 12'b111011101110;
20'b00110001100101111101: color_data = 12'b111011101110;
20'b00110001100101111110: color_data = 12'b111011101110;
20'b00110001100110000000: color_data = 12'b111011101110;
20'b00110001100110000001: color_data = 12'b111111111111;
20'b00110001100110000010: color_data = 12'b111011101110;
20'b00110001100110000011: color_data = 12'b111011101110;
20'b00110001100110000100: color_data = 12'b111011101110;
20'b00110001100110000110: color_data = 12'b111011101110;
20'b00110001100110000111: color_data = 12'b111011101110;
20'b00110001100110001000: color_data = 12'b111011101110;
20'b00110001100110001001: color_data = 12'b111111111111;
20'b00110001110011101011: color_data = 12'b111011101110;
20'b00110001110011101100: color_data = 12'b111011101110;
20'b00110001110011101101: color_data = 12'b111011101110;
20'b00110001110011101110: color_data = 12'b111011101110;
20'b00110001110011101111: color_data = 12'b111011101110;
20'b00110001110011110001: color_data = 12'b111011101110;
20'b00110001110011110010: color_data = 12'b111011101110;
20'b00110001110011110011: color_data = 12'b111011101110;
20'b00110001110011110100: color_data = 12'b111011101110;
20'b00110001110011110101: color_data = 12'b111011101110;
20'b00110001110100010111: color_data = 12'b111011101110;
20'b00110001110100011000: color_data = 12'b111011101110;
20'b00110001110100011001: color_data = 12'b111011101110;
20'b00110001110100011010: color_data = 12'b111011101110;
20'b00110001110100011011: color_data = 12'b111011101110;
20'b00110001110100011101: color_data = 12'b111011101110;
20'b00110001110100011110: color_data = 12'b111011101110;
20'b00110001110100011111: color_data = 12'b111011101110;
20'b00110001110100100000: color_data = 12'b111011101110;
20'b00110001110100100001: color_data = 12'b111011101110;
20'b00110001110100110011: color_data = 12'b111011101110;
20'b00110001110100110100: color_data = 12'b111011101110;
20'b00110001110100110101: color_data = 12'b111011101110;
20'b00110001110100110110: color_data = 12'b111011101110;
20'b00110001110100110111: color_data = 12'b111011101110;
20'b00110001110100111001: color_data = 12'b111011101110;
20'b00110001110100111010: color_data = 12'b111011101110;
20'b00110001110100111011: color_data = 12'b111011101110;
20'b00110001110100111100: color_data = 12'b111011101110;
20'b00110001110101000011: color_data = 12'b111011101110;
20'b00110001110101000100: color_data = 12'b111011101110;
20'b00110001110101000101: color_data = 12'b111011101110;
20'b00110001110101000110: color_data = 12'b111011101110;
20'b00110001110101000111: color_data = 12'b111011101110;
20'b00110001110101001001: color_data = 12'b111011101110;
20'b00110001110101001010: color_data = 12'b111011101110;
20'b00110001110101001011: color_data = 12'b111011101110;
20'b00110001110101001100: color_data = 12'b111011101110;
20'b00110001110101001101: color_data = 12'b111011101110;
20'b00110001110101010100: color_data = 12'b111011101110;
20'b00110001110101010101: color_data = 12'b111011101110;
20'b00110001110101010110: color_data = 12'b111011101110;
20'b00110001110101010111: color_data = 12'b111011101110;
20'b00110001110101011111: color_data = 12'b111011101110;
20'b00110001110101100000: color_data = 12'b111011101110;
20'b00110001110101100001: color_data = 12'b111011101110;
20'b00110001110101100010: color_data = 12'b111011101110;
20'b00110001110101100100: color_data = 12'b111011101110;
20'b00110001110101100101: color_data = 12'b111011101110;
20'b00110001110101100110: color_data = 12'b111011101110;
20'b00110001110101100111: color_data = 12'b111011101110;
20'b00110001110101101000: color_data = 12'b111011101110;
20'b00110001110101101111: color_data = 12'b111011101110;
20'b00110001110101110000: color_data = 12'b111011101110;
20'b00110001110101110001: color_data = 12'b111111111111;
20'b00110001110101110010: color_data = 12'b111011101110;
20'b00110001110101110011: color_data = 12'b111011101110;
20'b00110001110101110101: color_data = 12'b111011101110;
20'b00110001110101110110: color_data = 12'b111011101110;
20'b00110001110101110111: color_data = 12'b111011101110;
20'b00110001110101111000: color_data = 12'b111011101110;
20'b00110001110101111001: color_data = 12'b111111111111;
20'b00110001110101111011: color_data = 12'b111011101110;
20'b00110001110101111100: color_data = 12'b111111111111;
20'b00110001110101111101: color_data = 12'b111011101110;
20'b00110001110101111110: color_data = 12'b111111111111;
20'b00110001110110000000: color_data = 12'b111011101110;
20'b00110001110110000001: color_data = 12'b111011101110;
20'b00110001110110000010: color_data = 12'b111011101110;
20'b00110001110110000011: color_data = 12'b111011101110;
20'b00110001110110000100: color_data = 12'b111011101110;
20'b00110001110110000110: color_data = 12'b111011101110;
20'b00110001110110000111: color_data = 12'b111011101110;
20'b00110001110110001000: color_data = 12'b111011101110;
20'b00110001110110001001: color_data = 12'b111011101110;
20'b00110010000011101011: color_data = 12'b111011101110;
20'b00110010000011101100: color_data = 12'b111011101110;
20'b00110010000011101101: color_data = 12'b111011101110;
20'b00110010000011101110: color_data = 12'b111011101110;
20'b00110010000011101111: color_data = 12'b111011101110;
20'b00110010000011110001: color_data = 12'b111011101110;
20'b00110010000011110010: color_data = 12'b111011101110;
20'b00110010000011110011: color_data = 12'b111011101110;
20'b00110010000011110100: color_data = 12'b111011101110;
20'b00110010000011110101: color_data = 12'b111011101110;
20'b00110010000100010111: color_data = 12'b111011101110;
20'b00110010000100011000: color_data = 12'b111011101110;
20'b00110010000100011001: color_data = 12'b111011101110;
20'b00110010000100011010: color_data = 12'b111111111111;
20'b00110010000100011011: color_data = 12'b111011101110;
20'b00110010000100011101: color_data = 12'b111011101110;
20'b00110010000100011110: color_data = 12'b111011101110;
20'b00110010000100011111: color_data = 12'b111011101110;
20'b00110010000100100000: color_data = 12'b111011101110;
20'b00110010000100100001: color_data = 12'b111011101110;
20'b00110010000100110011: color_data = 12'b111011101110;
20'b00110010000100110100: color_data = 12'b111011101110;
20'b00110010000100110101: color_data = 12'b111011101110;
20'b00110010000100110110: color_data = 12'b111011101110;
20'b00110010000100110111: color_data = 12'b111011101110;
20'b00110010000100111001: color_data = 12'b111011101110;
20'b00110010000100111010: color_data = 12'b111011101110;
20'b00110010000100111011: color_data = 12'b111011101110;
20'b00110010000100111100: color_data = 12'b111011101110;
20'b00110010000101000011: color_data = 12'b111011101110;
20'b00110010000101000100: color_data = 12'b111011101110;
20'b00110010000101000101: color_data = 12'b111011101110;
20'b00110010000101000110: color_data = 12'b111011101110;
20'b00110010000101000111: color_data = 12'b111011101110;
20'b00110010000101001001: color_data = 12'b111011101110;
20'b00110010000101001010: color_data = 12'b111011101110;
20'b00110010000101001011: color_data = 12'b111011101110;
20'b00110010000101001100: color_data = 12'b111011101110;
20'b00110010000101001101: color_data = 12'b111011101110;
20'b00110010000101010100: color_data = 12'b111011101110;
20'b00110010000101010101: color_data = 12'b111011101110;
20'b00110010000101010110: color_data = 12'b111011101110;
20'b00110010000101010111: color_data = 12'b111011101110;
20'b00110010000101011111: color_data = 12'b111011101110;
20'b00110010000101100000: color_data = 12'b111011101110;
20'b00110010000101100001: color_data = 12'b111011101110;
20'b00110010000101100010: color_data = 12'b111011101110;
20'b00110010000101100100: color_data = 12'b111011101110;
20'b00110010000101100101: color_data = 12'b111011101110;
20'b00110010000101100110: color_data = 12'b111011101110;
20'b00110010000101100111: color_data = 12'b111011101110;
20'b00110010000101101000: color_data = 12'b111011101110;
20'b00110010000101101111: color_data = 12'b111011101110;
20'b00110010000101110000: color_data = 12'b111011101110;
20'b00110010000101110001: color_data = 12'b111011101110;
20'b00110010000101110010: color_data = 12'b111011101110;
20'b00110010000101110011: color_data = 12'b111011101110;
20'b00110010000101110101: color_data = 12'b111011101110;
20'b00110010000101110110: color_data = 12'b111011101110;
20'b00110010000101110111: color_data = 12'b111011101110;
20'b00110010000101111000: color_data = 12'b111011101110;
20'b00110010000101111001: color_data = 12'b111111111111;
20'b00110010000101111011: color_data = 12'b111011101110;
20'b00110010000101111100: color_data = 12'b111111111111;
20'b00110010000101111101: color_data = 12'b111011101110;
20'b00110010000101111110: color_data = 12'b111111111111;
20'b00110010000110000000: color_data = 12'b111011101110;
20'b00110010000110000001: color_data = 12'b111011101110;
20'b00110010000110000010: color_data = 12'b111011101110;
20'b00110010000110000011: color_data = 12'b111011101110;
20'b00110010000110000100: color_data = 12'b111011101110;
20'b00110010000110000110: color_data = 12'b111011101110;
20'b00110010000110000111: color_data = 12'b111011101110;
20'b00110010000110001000: color_data = 12'b111011101110;
20'b00110010000110001001: color_data = 12'b111011101110;
20'b00110010010011101011: color_data = 12'b111011101110;
20'b00110010010011101100: color_data = 12'b111011101110;
20'b00110010010011101101: color_data = 12'b111011101110;
20'b00110010010011101110: color_data = 12'b111111111111;
20'b00110010010011101111: color_data = 12'b111011101110;
20'b00110010010011110001: color_data = 12'b111011101110;
20'b00110010010011110010: color_data = 12'b111011101110;
20'b00110010010011110011: color_data = 12'b111011101110;
20'b00110010010011110100: color_data = 12'b111011101110;
20'b00110010010011110101: color_data = 12'b111011101110;
20'b00110010010100010111: color_data = 12'b111011101110;
20'b00110010010100011000: color_data = 12'b111011101110;
20'b00110010010100011001: color_data = 12'b111011101110;
20'b00110010010100011010: color_data = 12'b111011101110;
20'b00110010010100011011: color_data = 12'b111011101110;
20'b00110010010100011101: color_data = 12'b111011101110;
20'b00110010010100011110: color_data = 12'b111011101110;
20'b00110010010100011111: color_data = 12'b111011101110;
20'b00110010010100100000: color_data = 12'b111011101110;
20'b00110010010100100001: color_data = 12'b111011101110;
20'b00110010010100110011: color_data = 12'b111011101110;
20'b00110010010100110100: color_data = 12'b111111111111;
20'b00110010010100110101: color_data = 12'b111011101110;
20'b00110010010100110110: color_data = 12'b111011101110;
20'b00110010010100110111: color_data = 12'b111011101110;
20'b00110010010100111001: color_data = 12'b111011101110;
20'b00110010010100111010: color_data = 12'b111111111111;
20'b00110010010100111011: color_data = 12'b111011101110;
20'b00110010010100111100: color_data = 12'b111011101110;
20'b00110010010101000011: color_data = 12'b111011101110;
20'b00110010010101000100: color_data = 12'b111011101110;
20'b00110010010101000101: color_data = 12'b111011101110;
20'b00110010010101000110: color_data = 12'b111111111111;
20'b00110010010101000111: color_data = 12'b111011101110;
20'b00110010010101001001: color_data = 12'b111011101110;
20'b00110010010101001010: color_data = 12'b111011101110;
20'b00110010010101001011: color_data = 12'b111011101110;
20'b00110010010101001100: color_data = 12'b111011101110;
20'b00110010010101001101: color_data = 12'b111011101110;
20'b00110010010101010100: color_data = 12'b111011101110;
20'b00110010010101010101: color_data = 12'b111011101110;
20'b00110010010101010110: color_data = 12'b111011101110;
20'b00110010010101010111: color_data = 12'b111011101110;
20'b00110010010101011111: color_data = 12'b111011101110;
20'b00110010010101100000: color_data = 12'b111111111111;
20'b00110010010101100001: color_data = 12'b111011101110;
20'b00110010010101100010: color_data = 12'b111111111111;
20'b00110010010101100100: color_data = 12'b111011101110;
20'b00110010010101100101: color_data = 12'b111011101110;
20'b00110010010101100110: color_data = 12'b111011101110;
20'b00110010010101100111: color_data = 12'b111011101110;
20'b00110010010101101000: color_data = 12'b111011101110;
20'b00110010010101101111: color_data = 12'b111011101110;
20'b00110010010101110000: color_data = 12'b111011101110;
20'b00110010010101110001: color_data = 12'b111011101110;
20'b00110010010101110010: color_data = 12'b111011101110;
20'b00110010010101110011: color_data = 12'b111011101110;
20'b00110010010101110101: color_data = 12'b111111111111;
20'b00110010010101110110: color_data = 12'b111011101110;
20'b00110010010101110111: color_data = 12'b111111111111;
20'b00110010010101111000: color_data = 12'b111111111111;
20'b00110010010101111001: color_data = 12'b111011101110;
20'b00110010010101111011: color_data = 12'b111011101110;
20'b00110010010101111100: color_data = 12'b111011101110;
20'b00110010010101111101: color_data = 12'b111011101110;
20'b00110010010101111110: color_data = 12'b111011101110;
20'b00110010010110000000: color_data = 12'b111011101110;
20'b00110010010110000001: color_data = 12'b111111111111;
20'b00110010010110000010: color_data = 12'b111011101110;
20'b00110010010110000011: color_data = 12'b111011101110;
20'b00110010010110000100: color_data = 12'b111011101110;
20'b00110010010110000110: color_data = 12'b111011101110;
20'b00110010010110000111: color_data = 12'b111011101110;
20'b00110010010110001000: color_data = 12'b111011101110;
20'b00110010010110001001: color_data = 12'b111111111111;
20'b00110010100100000001: color_data = 12'b111111111111;
20'b00110010100100000010: color_data = 12'b111011101110;
20'b00110010100100000011: color_data = 12'b111011101110;
20'b00110010100100000100: color_data = 12'b111011101110;
20'b00110010100100000101: color_data = 12'b111011101110;
20'b00110010100100000111: color_data = 12'b111011101110;
20'b00110010100100001000: color_data = 12'b111011101110;
20'b00110010100100001001: color_data = 12'b111011101110;
20'b00110010100100001010: color_data = 12'b111011101110;
20'b00110010100100001011: color_data = 12'b111011101110;
20'b00110010100100001101: color_data = 12'b111111111111;
20'b00110010100100001110: color_data = 12'b111011101110;
20'b00110010100100001111: color_data = 12'b111111111111;
20'b00110010100100010000: color_data = 12'b111011101110;
20'b00110010100101010100: color_data = 12'b111011101110;
20'b00110010100101010101: color_data = 12'b111011101110;
20'b00110010100101010110: color_data = 12'b111011101110;
20'b00110010100101010111: color_data = 12'b111011101110;
20'b00110010110011101011: color_data = 12'b111011101110;
20'b00110010110011101100: color_data = 12'b111011101110;
20'b00110010110011101101: color_data = 12'b111111111111;
20'b00110010110011101110: color_data = 12'b111011101110;
20'b00110010110011101111: color_data = 12'b111011101110;
20'b00110010110011110001: color_data = 12'b111011101110;
20'b00110010110011110010: color_data = 12'b111011101110;
20'b00110010110011110011: color_data = 12'b111011101110;
20'b00110010110011110100: color_data = 12'b111011101110;
20'b00110010110011110101: color_data = 12'b111011101110;
20'b00110010110100000001: color_data = 12'b111011101110;
20'b00110010110100000010: color_data = 12'b111011101110;
20'b00110010110100000011: color_data = 12'b111011101110;
20'b00110010110100000100: color_data = 12'b111011101110;
20'b00110010110100000101: color_data = 12'b111011101110;
20'b00110010110100000111: color_data = 12'b111011101110;
20'b00110010110100001000: color_data = 12'b111011101110;
20'b00110010110100001001: color_data = 12'b111011101110;
20'b00110010110100001010: color_data = 12'b111011101110;
20'b00110010110100001011: color_data = 12'b111011101110;
20'b00110010110100001101: color_data = 12'b111011101110;
20'b00110010110100001110: color_data = 12'b111011101110;
20'b00110010110100001111: color_data = 12'b111011101110;
20'b00110010110100010000: color_data = 12'b111111111111;
20'b00110010110100010111: color_data = 12'b111011101110;
20'b00110010110100011000: color_data = 12'b111011101110;
20'b00110010110100011001: color_data = 12'b111011101110;
20'b00110010110100011010: color_data = 12'b111011101110;
20'b00110010110100011011: color_data = 12'b111011101110;
20'b00110010110100011101: color_data = 12'b111011101110;
20'b00110010110100011110: color_data = 12'b111011101110;
20'b00110010110100011111: color_data = 12'b111011101110;
20'b00110010110100100000: color_data = 12'b111011101110;
20'b00110010110100100001: color_data = 12'b111011101110;
20'b00110010110100100011: color_data = 12'b111011101110;
20'b00110010110100100100: color_data = 12'b111011101110;
20'b00110010110100100101: color_data = 12'b111011101110;
20'b00110010110100100110: color_data = 12'b111011101110;
20'b00110010110100101000: color_data = 12'b111011101110;
20'b00110010110100101001: color_data = 12'b111111111111;
20'b00110010110100101010: color_data = 12'b111011101110;
20'b00110010110100101011: color_data = 12'b111011101110;
20'b00110010110100101100: color_data = 12'b111011101110;
20'b00110010110100101110: color_data = 12'b111011101110;
20'b00110010110100101111: color_data = 12'b111111111111;
20'b00110010110100110000: color_data = 12'b111011101110;
20'b00110010110100110001: color_data = 12'b111011101110;
20'b00110010110100110011: color_data = 12'b111111111111;
20'b00110010110100110100: color_data = 12'b111011101110;
20'b00110010110100110101: color_data = 12'b111011101110;
20'b00110010110100110110: color_data = 12'b111011101110;
20'b00110010110100110111: color_data = 12'b111011101110;
20'b00110010110100111001: color_data = 12'b111011101110;
20'b00110010110100111010: color_data = 12'b111111111111;
20'b00110010110100111011: color_data = 12'b111111111111;
20'b00110010110100111100: color_data = 12'b111011101110;
20'b00110010110101000011: color_data = 12'b111011101110;
20'b00110010110101000100: color_data = 12'b111011101110;
20'b00110010110101000101: color_data = 12'b111111111111;
20'b00110010110101000110: color_data = 12'b111011101110;
20'b00110010110101000111: color_data = 12'b111011101110;
20'b00110010110101001001: color_data = 12'b111011101110;
20'b00110010110101001010: color_data = 12'b111011101110;
20'b00110010110101001011: color_data = 12'b111011101110;
20'b00110010110101001100: color_data = 12'b111011101110;
20'b00110010110101001101: color_data = 12'b111011101110;
20'b00110010110101011111: color_data = 12'b111011101110;
20'b00110010110101100000: color_data = 12'b111011101110;
20'b00110010110101100001: color_data = 12'b111011101110;
20'b00110010110101100010: color_data = 12'b111011101110;
20'b00110010110101100100: color_data = 12'b111011101110;
20'b00110010110101100101: color_data = 12'b111011101110;
20'b00110010110101100110: color_data = 12'b111011101110;
20'b00110010110101100111: color_data = 12'b111011101110;
20'b00110010110101101000: color_data = 12'b111011101110;
20'b00110010110101101111: color_data = 12'b111011101110;
20'b00110010110101110000: color_data = 12'b111011101110;
20'b00110010110101110001: color_data = 12'b111011101110;
20'b00110010110101110010: color_data = 12'b111011101110;
20'b00110010110101110011: color_data = 12'b111011101110;
20'b00110010110101110101: color_data = 12'b111011101110;
20'b00110010110101110110: color_data = 12'b111011101110;
20'b00110010110101110111: color_data = 12'b111011101110;
20'b00110010110101111000: color_data = 12'b111011101110;
20'b00110010110101111001: color_data = 12'b111011101110;
20'b00110011000011101011: color_data = 12'b111111111111;
20'b00110011000011101100: color_data = 12'b111011101110;
20'b00110011000011101101: color_data = 12'b111011101110;
20'b00110011000011101110: color_data = 12'b111011101110;
20'b00110011000011101111: color_data = 12'b111011101110;
20'b00110011000011110001: color_data = 12'b111011101110;
20'b00110011000011110010: color_data = 12'b111111111111;
20'b00110011000011110011: color_data = 12'b111011101110;
20'b00110011000011110100: color_data = 12'b111011101110;
20'b00110011000011110101: color_data = 12'b111011101110;
20'b00110011000100000001: color_data = 12'b111011101110;
20'b00110011000100000010: color_data = 12'b111011101110;
20'b00110011000100000011: color_data = 12'b111111111111;
20'b00110011000100000100: color_data = 12'b111011101110;
20'b00110011000100000101: color_data = 12'b111011101110;
20'b00110011000100000111: color_data = 12'b111011101110;
20'b00110011000100001000: color_data = 12'b111011101110;
20'b00110011000100001001: color_data = 12'b111011101110;
20'b00110011000100001010: color_data = 12'b111111111111;
20'b00110011000100001011: color_data = 12'b111011101110;
20'b00110011000100001101: color_data = 12'b111011101110;
20'b00110011000100001110: color_data = 12'b111011101110;
20'b00110011000100001111: color_data = 12'b111011101110;
20'b00110011000100010000: color_data = 12'b111011101110;
20'b00110011000100010111: color_data = 12'b111011101110;
20'b00110011000100011000: color_data = 12'b111011101110;
20'b00110011000100011001: color_data = 12'b111011101110;
20'b00110011000100011010: color_data = 12'b111011101110;
20'b00110011000100011011: color_data = 12'b111011101110;
20'b00110011000100011101: color_data = 12'b111111111111;
20'b00110011000100011110: color_data = 12'b111011101110;
20'b00110011000100011111: color_data = 12'b111011101110;
20'b00110011000100100000: color_data = 12'b111011101110;
20'b00110011000100100001: color_data = 12'b111011101110;
20'b00110011000100100011: color_data = 12'b111111111111;
20'b00110011000100100100: color_data = 12'b111011101110;
20'b00110011000100100101: color_data = 12'b111011101110;
20'b00110011000100100110: color_data = 12'b111011101110;
20'b00110011000100101000: color_data = 12'b111011101110;
20'b00110011000100101001: color_data = 12'b111011101110;
20'b00110011000100101010: color_data = 12'b111111111111;
20'b00110011000100101011: color_data = 12'b111011101110;
20'b00110011000100101100: color_data = 12'b111011101110;
20'b00110011000100101110: color_data = 12'b111011101110;
20'b00110011000100101111: color_data = 12'b111011101110;
20'b00110011000100110000: color_data = 12'b111011101110;
20'b00110011000100110001: color_data = 12'b111011101110;
20'b00110011000100110011: color_data = 12'b111011101110;
20'b00110011000100110100: color_data = 12'b111011101110;
20'b00110011000100110101: color_data = 12'b111011101110;
20'b00110011000100110110: color_data = 12'b111011101110;
20'b00110011000100110111: color_data = 12'b111011101110;
20'b00110011000100111001: color_data = 12'b111011101110;
20'b00110011000100111010: color_data = 12'b111011101110;
20'b00110011000100111011: color_data = 12'b111011101110;
20'b00110011000100111100: color_data = 12'b111011101110;
20'b00110011000101000011: color_data = 12'b111111111111;
20'b00110011000101000100: color_data = 12'b111011101110;
20'b00110011000101000101: color_data = 12'b111011101110;
20'b00110011000101000110: color_data = 12'b111011101110;
20'b00110011000101000111: color_data = 12'b111011101110;
20'b00110011000101001001: color_data = 12'b111011101110;
20'b00110011000101001010: color_data = 12'b111111111111;
20'b00110011000101001011: color_data = 12'b111011101110;
20'b00110011000101001100: color_data = 12'b111011101110;
20'b00110011000101001101: color_data = 12'b111011101110;
20'b00110011000101011111: color_data = 12'b111111111111;
20'b00110011000101100000: color_data = 12'b111011101110;
20'b00110011000101100001: color_data = 12'b111011101110;
20'b00110011000101100010: color_data = 12'b111011101110;
20'b00110011000101100100: color_data = 12'b111011101110;
20'b00110011000101100101: color_data = 12'b111111111111;
20'b00110011000101100110: color_data = 12'b111111111111;
20'b00110011000101100111: color_data = 12'b111011101110;
20'b00110011000101101000: color_data = 12'b111011101110;
20'b00110011000101101111: color_data = 12'b111011101110;
20'b00110011000101110000: color_data = 12'b111011101110;
20'b00110011000101110001: color_data = 12'b111111111111;
20'b00110011000101110010: color_data = 12'b111111111111;
20'b00110011000101110011: color_data = 12'b111011101110;
20'b00110011000101110101: color_data = 12'b111011101110;
20'b00110011000101110110: color_data = 12'b111011101110;
20'b00110011000101110111: color_data = 12'b111011101110;
20'b00110011000101111000: color_data = 12'b111011101110;
20'b00110011000101111001: color_data = 12'b111011101110;
20'b00110011010011101011: color_data = 12'b111011101110;
20'b00110011010011101100: color_data = 12'b111011101110;
20'b00110011010011101101: color_data = 12'b111011101110;
20'b00110011010011101110: color_data = 12'b111011101110;
20'b00110011010011101111: color_data = 12'b111011101110;
20'b00110011010011110001: color_data = 12'b111011101110;
20'b00110011010011110010: color_data = 12'b111011101110;
20'b00110011010011110011: color_data = 12'b111111111111;
20'b00110011010011110100: color_data = 12'b111111111111;
20'b00110011010011110101: color_data = 12'b111011101110;
20'b00110011010100000001: color_data = 12'b111011101110;
20'b00110011010100000010: color_data = 12'b111011101110;
20'b00110011010100000011: color_data = 12'b111011101110;
20'b00110011010100000100: color_data = 12'b111011101110;
20'b00110011010100000101: color_data = 12'b111011101110;
20'b00110011010100000111: color_data = 12'b111011101110;
20'b00110011010100001000: color_data = 12'b111011101110;
20'b00110011010100001001: color_data = 12'b111111111111;
20'b00110011010100001010: color_data = 12'b111011101110;
20'b00110011010100001011: color_data = 12'b111011101110;
20'b00110011010100001101: color_data = 12'b111011101110;
20'b00110011010100001110: color_data = 12'b111011101110;
20'b00110011010100001111: color_data = 12'b111011101110;
20'b00110011010100010000: color_data = 12'b111111111111;
20'b00110011010100010111: color_data = 12'b111011101110;
20'b00110011010100011000: color_data = 12'b111011101110;
20'b00110011010100011001: color_data = 12'b111011101110;
20'b00110011010100011010: color_data = 12'b111011101110;
20'b00110011010100011011: color_data = 12'b111111111111;
20'b00110011010100011101: color_data = 12'b111011101110;
20'b00110011010100011110: color_data = 12'b111011101110;
20'b00110011010100011111: color_data = 12'b111011101110;
20'b00110011010100100000: color_data = 12'b111011101110;
20'b00110011010100100001: color_data = 12'b111111111111;
20'b00110011010100100011: color_data = 12'b111011101110;
20'b00110011010100100100: color_data = 12'b111011101110;
20'b00110011010100100101: color_data = 12'b111011101110;
20'b00110011010100100110: color_data = 12'b111011101110;
20'b00110011010100101000: color_data = 12'b111011101110;
20'b00110011010100101001: color_data = 12'b111011101110;
20'b00110011010100101010: color_data = 12'b111011101110;
20'b00110011010100101011: color_data = 12'b111011101110;
20'b00110011010100101100: color_data = 12'b111011101110;
20'b00110011010100101110: color_data = 12'b111011101110;
20'b00110011010100101111: color_data = 12'b111011101110;
20'b00110011010100110000: color_data = 12'b111011101110;
20'b00110011010100110001: color_data = 12'b111111111111;
20'b00110011010100110011: color_data = 12'b111011101110;
20'b00110011010100110100: color_data = 12'b111111111111;
20'b00110011010100110101: color_data = 12'b111011101110;
20'b00110011010100110110: color_data = 12'b111011101110;
20'b00110011010100110111: color_data = 12'b111011101110;
20'b00110011010100111001: color_data = 12'b111011101110;
20'b00110011010100111010: color_data = 12'b111111111111;
20'b00110011010100111011: color_data = 12'b111011101110;
20'b00110011010100111100: color_data = 12'b111011101110;
20'b00110011010101000011: color_data = 12'b111011101110;
20'b00110011010101000100: color_data = 12'b111011101110;
20'b00110011010101000101: color_data = 12'b111011101110;
20'b00110011010101000110: color_data = 12'b111011101110;
20'b00110011010101000111: color_data = 12'b111011101110;
20'b00110011010101001001: color_data = 12'b111011101110;
20'b00110011010101001010: color_data = 12'b111011101110;
20'b00110011010101001011: color_data = 12'b111111111111;
20'b00110011010101001100: color_data = 12'b111111111111;
20'b00110011010101001101: color_data = 12'b111011101110;
20'b00110011010101011111: color_data = 12'b111011101110;
20'b00110011010101100000: color_data = 12'b111011101110;
20'b00110011010101100001: color_data = 12'b111111111111;
20'b00110011010101100010: color_data = 12'b111011101110;
20'b00110011010101100100: color_data = 12'b111011101110;
20'b00110011010101100101: color_data = 12'b111011101110;
20'b00110011010101100110: color_data = 12'b111011101110;
20'b00110011010101100111: color_data = 12'b111011101110;
20'b00110011010101101000: color_data = 12'b111011101110;
20'b00110011010101101111: color_data = 12'b111011101110;
20'b00110011010101110000: color_data = 12'b111011101110;
20'b00110011010101110001: color_data = 12'b111011101110;
20'b00110011010101110010: color_data = 12'b111011101110;
20'b00110011010101110011: color_data = 12'b111011101110;
20'b00110011010101110101: color_data = 12'b111011101110;
20'b00110011010101110110: color_data = 12'b111111111111;
20'b00110011010101110111: color_data = 12'b111011101110;
20'b00110011010101111000: color_data = 12'b111011101110;
20'b00110011010101111001: color_data = 12'b111011101110;
20'b00110011100011101011: color_data = 12'b111011101110;
20'b00110011100011101100: color_data = 12'b111011101110;
20'b00110011100011101101: color_data = 12'b111011101110;
20'b00110011100011101110: color_data = 12'b111011101110;
20'b00110011100011101111: color_data = 12'b111011101110;
20'b00110011100011110001: color_data = 12'b111011101110;
20'b00110011100011110010: color_data = 12'b111011101110;
20'b00110011100011110011: color_data = 12'b111011101110;
20'b00110011100011110100: color_data = 12'b111011101110;
20'b00110011100011110101: color_data = 12'b111111111111;
20'b00110011100100000001: color_data = 12'b111011101110;
20'b00110011100100000010: color_data = 12'b111011101110;
20'b00110011100100000011: color_data = 12'b111111111111;
20'b00110011100100000100: color_data = 12'b111011101110;
20'b00110011100100000101: color_data = 12'b111111111111;
20'b00110011100100000111: color_data = 12'b111011101110;
20'b00110011100100001000: color_data = 12'b111011101110;
20'b00110011100100001001: color_data = 12'b111011101110;
20'b00110011100100001010: color_data = 12'b111111111111;
20'b00110011100100001011: color_data = 12'b111011101110;
20'b00110011100100001101: color_data = 12'b111011101110;
20'b00110011100100001110: color_data = 12'b111111111111;
20'b00110011100100001111: color_data = 12'b111011101110;
20'b00110011100100010000: color_data = 12'b111011101110;
20'b00110011100100010111: color_data = 12'b111011101110;
20'b00110011100100011000: color_data = 12'b111011101110;
20'b00110011100100011001: color_data = 12'b111011101110;
20'b00110011100100011010: color_data = 12'b111011101110;
20'b00110011100100011011: color_data = 12'b111011101110;
20'b00110011100100011101: color_data = 12'b111111111111;
20'b00110011100100011110: color_data = 12'b111011101110;
20'b00110011100100011111: color_data = 12'b111111111111;
20'b00110011100100100000: color_data = 12'b111111111111;
20'b00110011100100100001: color_data = 12'b111011101110;
20'b00110011100100100011: color_data = 12'b111111111111;
20'b00110011100100100100: color_data = 12'b111011101110;
20'b00110011100100100101: color_data = 12'b111111111111;
20'b00110011100100100110: color_data = 12'b111011101110;
20'b00110011100100101000: color_data = 12'b111011101110;
20'b00110011100100101001: color_data = 12'b111011101110;
20'b00110011100100101010: color_data = 12'b111011101110;
20'b00110011100100101011: color_data = 12'b111011101110;
20'b00110011100100101100: color_data = 12'b111011101110;
20'b00110011100100101110: color_data = 12'b111011101110;
20'b00110011100100101111: color_data = 12'b111011101110;
20'b00110011100100110000: color_data = 12'b111011101110;
20'b00110011100100110001: color_data = 12'b111111111111;
20'b00110011100100110011: color_data = 12'b111011101110;
20'b00110011100100110100: color_data = 12'b111011101110;
20'b00110011100100110101: color_data = 12'b111011101110;
20'b00110011100100110110: color_data = 12'b111011101110;
20'b00110011100100110111: color_data = 12'b111011101110;
20'b00110011100100111001: color_data = 12'b111011101110;
20'b00110011100100111010: color_data = 12'b111011101110;
20'b00110011100100111011: color_data = 12'b111011101110;
20'b00110011100100111100: color_data = 12'b111011101110;
20'b00110011100101000011: color_data = 12'b111011101110;
20'b00110011100101000100: color_data = 12'b111011101110;
20'b00110011100101000101: color_data = 12'b111011101110;
20'b00110011100101000110: color_data = 12'b111011101110;
20'b00110011100101000111: color_data = 12'b111011101110;
20'b00110011100101001001: color_data = 12'b111011101110;
20'b00110011100101001010: color_data = 12'b111011101110;
20'b00110011100101001011: color_data = 12'b111011101110;
20'b00110011100101001100: color_data = 12'b111011101110;
20'b00110011100101001101: color_data = 12'b111111111111;
20'b00110011100101011111: color_data = 12'b111011101110;
20'b00110011100101100000: color_data = 12'b111011101110;
20'b00110011100101100001: color_data = 12'b111011101110;
20'b00110011100101100010: color_data = 12'b111011101110;
20'b00110011100101100100: color_data = 12'b111011101110;
20'b00110011100101100101: color_data = 12'b111011101110;
20'b00110011100101100110: color_data = 12'b111111111111;
20'b00110011100101100111: color_data = 12'b111111111111;
20'b00110011100101101000: color_data = 12'b111011101110;
20'b00110011100101101111: color_data = 12'b111011101110;
20'b00110011100101110000: color_data = 12'b111111111111;
20'b00110011100101110001: color_data = 12'b111111111111;
20'b00110011100101110010: color_data = 12'b111011101110;
20'b00110011100101110011: color_data = 12'b111011101110;
20'b00110011100101110101: color_data = 12'b111011101110;
20'b00110011100101110110: color_data = 12'b111011101110;
20'b00110011100101110111: color_data = 12'b111011101110;
20'b00110011100101111000: color_data = 12'b111011101110;
20'b00110011100101111001: color_data = 12'b111011101110;
20'b00110011110100010111: color_data = 12'b111011101110;
20'b00110011110100011000: color_data = 12'b111011101110;
20'b00110011110100011001: color_data = 12'b111011101110;
20'b00110011110100011010: color_data = 12'b111011101110;
20'b00110011110100011011: color_data = 12'b111011101110;
20'b00110011110100011101: color_data = 12'b111011101110;
20'b00110011110100011110: color_data = 12'b111111111111;
20'b00110011110100011111: color_data = 12'b111011101110;
20'b00110011110100100000: color_data = 12'b111011101110;
20'b00110011110100100001: color_data = 12'b111011101110;
20'b00110011110100100011: color_data = 12'b111011101110;
20'b00110011110100100100: color_data = 12'b111011101110;
20'b00110011110100100101: color_data = 12'b111011101110;
20'b00110011110100100110: color_data = 12'b111011101110;
20'b00110011110100101000: color_data = 12'b111011101110;
20'b00110011110100101001: color_data = 12'b111011101110;
20'b00110011110100101010: color_data = 12'b111011101110;
20'b00110011110100101011: color_data = 12'b111011101110;
20'b00110011110100101100: color_data = 12'b111011101110;
20'b00110011110100101110: color_data = 12'b111011101110;
20'b00110011110100101111: color_data = 12'b111011101110;
20'b00110011110100110000: color_data = 12'b111111111111;
20'b00110011110100110001: color_data = 12'b111011101110;
20'b00110011110100110011: color_data = 12'b111011101110;
20'b00110011110100110100: color_data = 12'b111011101110;
20'b00110011110100110101: color_data = 12'b111011101110;
20'b00110011110100110110: color_data = 12'b111011101110;
20'b00110011110100110111: color_data = 12'b111011101110;
20'b00110011110100111001: color_data = 12'b111111111111;
20'b00110011110100111010: color_data = 12'b111011101110;
20'b00110011110100111011: color_data = 12'b111011101110;
20'b00110011110100111100: color_data = 12'b111011101110;
20'b00110100000011101011: color_data = 12'b111011101110;
20'b00110100000011101100: color_data = 12'b111011101110;
20'b00110100000011101101: color_data = 12'b111111111111;
20'b00110100000011101110: color_data = 12'b111011101110;
20'b00110100000011101111: color_data = 12'b111011101110;
20'b00110100000011110001: color_data = 12'b111011101110;
20'b00110100000011110010: color_data = 12'b111011101110;
20'b00110100000011110011: color_data = 12'b111011101110;
20'b00110100000011110100: color_data = 12'b111011101110;
20'b00110100000011110101: color_data = 12'b111111111111;
20'b00110100000100000111: color_data = 12'b111011101110;
20'b00110100000100001000: color_data = 12'b111011101110;
20'b00110100000100001001: color_data = 12'b111011101110;
20'b00110100000100001010: color_data = 12'b111011101110;
20'b00110100000100001011: color_data = 12'b111011101110;
20'b00110100000100001101: color_data = 12'b111011101110;
20'b00110100000100001110: color_data = 12'b111011101110;
20'b00110100000100001111: color_data = 12'b111011101110;
20'b00110100000100010000: color_data = 12'b111111111111;
20'b00110100000101000011: color_data = 12'b111011101110;
20'b00110100000101000100: color_data = 12'b111011101110;
20'b00110100000101000101: color_data = 12'b111011101110;
20'b00110100000101000110: color_data = 12'b111011101110;
20'b00110100000101000111: color_data = 12'b111011101110;
20'b00110100000101001001: color_data = 12'b111011101110;
20'b00110100000101001010: color_data = 12'b111011101110;
20'b00110100000101001011: color_data = 12'b111011101110;
20'b00110100000101001100: color_data = 12'b111011101110;
20'b00110100000101001101: color_data = 12'b111011101110;
20'b00110100000101011111: color_data = 12'b111011101110;
20'b00110100000101100000: color_data = 12'b111011101110;
20'b00110100000101100001: color_data = 12'b111111111111;
20'b00110100000101100010: color_data = 12'b111011101110;
20'b00110100000101100100: color_data = 12'b111011101110;
20'b00110100000101100101: color_data = 12'b111011101110;
20'b00110100000101100110: color_data = 12'b111011101110;
20'b00110100000101100111: color_data = 12'b111011101110;
20'b00110100000101101000: color_data = 12'b111011101110;
20'b00110100000101101111: color_data = 12'b111011101110;
20'b00110100000101110000: color_data = 12'b111011101110;
20'b00110100000101110001: color_data = 12'b111011101110;
20'b00110100000101110010: color_data = 12'b111011101110;
20'b00110100000101110011: color_data = 12'b111011101110;
20'b00110100000101110101: color_data = 12'b111011101110;
20'b00110100000101110110: color_data = 12'b111111111111;
20'b00110100000101110111: color_data = 12'b111011101110;
20'b00110100000101111000: color_data = 12'b111111111111;
20'b00110100000101111001: color_data = 12'b111011101110;
20'b00110100010011101011: color_data = 12'b111011101110;
20'b00110100010011101100: color_data = 12'b111011101110;
20'b00110100010011101101: color_data = 12'b111011101110;
20'b00110100010011101110: color_data = 12'b111011101110;
20'b00110100010011101111: color_data = 12'b111011101110;
20'b00110100010011110001: color_data = 12'b111011101110;
20'b00110100010011110010: color_data = 12'b111011101110;
20'b00110100010011110011: color_data = 12'b111011101110;
20'b00110100010011110100: color_data = 12'b111011101110;
20'b00110100010011110101: color_data = 12'b111011101110;
20'b00110100010100000111: color_data = 12'b111011101110;
20'b00110100010100001000: color_data = 12'b111011101110;
20'b00110100010100001001: color_data = 12'b111011101110;
20'b00110100010100001010: color_data = 12'b111011101110;
20'b00110100010100001011: color_data = 12'b111111111111;
20'b00110100010100001101: color_data = 12'b111011101110;
20'b00110100010100001110: color_data = 12'b111011101110;
20'b00110100010100001111: color_data = 12'b111011101110;
20'b00110100010100010000: color_data = 12'b111011101110;
20'b00110100010100010111: color_data = 12'b111011101110;
20'b00110100010100011000: color_data = 12'b111111111111;
20'b00110100010100011001: color_data = 12'b111111111111;
20'b00110100010100011010: color_data = 12'b111011101110;
20'b00110100010100011011: color_data = 12'b111011101110;
20'b00110100010100011101: color_data = 12'b111011101110;
20'b00110100010100011110: color_data = 12'b111011101110;
20'b00110100010100011111: color_data = 12'b111011101110;
20'b00110100010100100000: color_data = 12'b111011101110;
20'b00110100010100100001: color_data = 12'b111111111111;
20'b00110100010100110011: color_data = 12'b111011101110;
20'b00110100010100110100: color_data = 12'b111011101110;
20'b00110100010100110101: color_data = 12'b111011101110;
20'b00110100010100110110: color_data = 12'b111011101110;
20'b00110100010100110111: color_data = 12'b111011101110;
20'b00110100010100111001: color_data = 12'b111011101110;
20'b00110100010100111010: color_data = 12'b111011101110;
20'b00110100010100111011: color_data = 12'b111011101110;
20'b00110100010100111100: color_data = 12'b111011101110;
20'b00110100010101000011: color_data = 12'b111111111111;
20'b00110100010101000100: color_data = 12'b111011101110;
20'b00110100010101000101: color_data = 12'b111111111111;
20'b00110100010101000110: color_data = 12'b111011101110;
20'b00110100010101000111: color_data = 12'b111011101110;
20'b00110100010101001001: color_data = 12'b111011101110;
20'b00110100010101001010: color_data = 12'b111011101110;
20'b00110100010101001011: color_data = 12'b111011101110;
20'b00110100010101001100: color_data = 12'b111011101110;
20'b00110100010101001101: color_data = 12'b111011101110;
20'b00110100010101011111: color_data = 12'b111011101110;
20'b00110100010101100000: color_data = 12'b111111111111;
20'b00110100010101100001: color_data = 12'b111011101110;
20'b00110100010101100010: color_data = 12'b111111111111;
20'b00110100010101100100: color_data = 12'b111011101110;
20'b00110100010101100101: color_data = 12'b111011101110;
20'b00110100010101100110: color_data = 12'b111011101110;
20'b00110100010101100111: color_data = 12'b111011101110;
20'b00110100010101101000: color_data = 12'b111011101110;
20'b00110100010101101111: color_data = 12'b111011101110;
20'b00110100010101110000: color_data = 12'b111011101110;
20'b00110100010101110001: color_data = 12'b111011101110;
20'b00110100010101110010: color_data = 12'b111011101110;
20'b00110100010101110011: color_data = 12'b111011101110;
20'b00110100010101110101: color_data = 12'b111111111111;
20'b00110100010101110110: color_data = 12'b111011101110;
20'b00110100010101110111: color_data = 12'b111111111111;
20'b00110100010101111000: color_data = 12'b111011101110;
20'b00110100010101111001: color_data = 12'b111111111111;
20'b00110100100011101011: color_data = 12'b111011101110;
20'b00110100100011101100: color_data = 12'b111011101110;
20'b00110100100011101101: color_data = 12'b111111111111;
20'b00110100100011101110: color_data = 12'b111011101110;
20'b00110100100011101111: color_data = 12'b111011101110;
20'b00110100100011110001: color_data = 12'b111011101110;
20'b00110100100011110010: color_data = 12'b111111111111;
20'b00110100100011110011: color_data = 12'b111011101110;
20'b00110100100011110100: color_data = 12'b111011101110;
20'b00110100100011110101: color_data = 12'b111011101110;
20'b00110100100100000111: color_data = 12'b111111111111;
20'b00110100100100001000: color_data = 12'b111011101110;
20'b00110100100100001001: color_data = 12'b111011101110;
20'b00110100100100001010: color_data = 12'b111111111111;
20'b00110100100100001011: color_data = 12'b111011101110;
20'b00110100100100001101: color_data = 12'b111011101110;
20'b00110100100100001110: color_data = 12'b111111111111;
20'b00110100100100001111: color_data = 12'b111011101110;
20'b00110100100100010000: color_data = 12'b111111111111;
20'b00110100100100010111: color_data = 12'b111011101110;
20'b00110100100100011000: color_data = 12'b111011101110;
20'b00110100100100011001: color_data = 12'b111011101110;
20'b00110100100100011010: color_data = 12'b111011101110;
20'b00110100100100011011: color_data = 12'b111011101110;
20'b00110100100100011101: color_data = 12'b111011101110;
20'b00110100100100011110: color_data = 12'b111111111111;
20'b00110100100100011111: color_data = 12'b111011101110;
20'b00110100100100100000: color_data = 12'b111011101110;
20'b00110100100100100001: color_data = 12'b111011101110;
20'b00110100100100110011: color_data = 12'b111011101110;
20'b00110100100100110100: color_data = 12'b111011101110;
20'b00110100100100110101: color_data = 12'b111011101110;
20'b00110100100100110110: color_data = 12'b111011101110;
20'b00110100100100110111: color_data = 12'b111011101110;
20'b00110100100100111001: color_data = 12'b111011101110;
20'b00110100100100111010: color_data = 12'b111011101110;
20'b00110100100100111011: color_data = 12'b111011101110;
20'b00110100100100111100: color_data = 12'b111111111111;
20'b00110100100101000011: color_data = 12'b111011101110;
20'b00110100100101000100: color_data = 12'b111111111111;
20'b00110100100101000101: color_data = 12'b111011101110;
20'b00110100100101000110: color_data = 12'b111011101110;
20'b00110100100101000111: color_data = 12'b111011101110;
20'b00110100100101001001: color_data = 12'b111011101110;
20'b00110100100101001010: color_data = 12'b111011101110;
20'b00110100100101001011: color_data = 12'b111011101110;
20'b00110100100101001100: color_data = 12'b111011101110;
20'b00110100100101001101: color_data = 12'b111011101110;
20'b00110100100101011111: color_data = 12'b111011101110;
20'b00110100100101100000: color_data = 12'b111011101110;
20'b00110100100101100001: color_data = 12'b111011101110;
20'b00110100100101100010: color_data = 12'b111011101110;
20'b00110100100101100100: color_data = 12'b111111111111;
20'b00110100100101100101: color_data = 12'b111011101110;
20'b00110100100101100110: color_data = 12'b111011101110;
20'b00110100100101100111: color_data = 12'b111011101110;
20'b00110100100101101000: color_data = 12'b111011101110;
20'b00110100100101101111: color_data = 12'b111011101110;
20'b00110100100101110000: color_data = 12'b111011101110;
20'b00110100100101110001: color_data = 12'b111011101110;
20'b00110100100101110010: color_data = 12'b111011101110;
20'b00110100100101110011: color_data = 12'b111111111111;
20'b00110100100101110101: color_data = 12'b111011101110;
20'b00110100100101110110: color_data = 12'b111011101110;
20'b00110100100101110111: color_data = 12'b111011101110;
20'b00110100100101111000: color_data = 12'b111111111111;
20'b00110100100101111001: color_data = 12'b111111111111;
20'b00110100110011101011: color_data = 12'b111111111111;
20'b00110100110011101100: color_data = 12'b111011101110;
20'b00110100110011101101: color_data = 12'b111011101110;
20'b00110100110011101110: color_data = 12'b111011101110;
20'b00110100110011101111: color_data = 12'b111011101110;
20'b00110100110011110001: color_data = 12'b111011101110;
20'b00110100110011110010: color_data = 12'b111011101110;
20'b00110100110011110011: color_data = 12'b111011101110;
20'b00110100110011110100: color_data = 12'b111111111111;
20'b00110100110011110101: color_data = 12'b111011101110;
20'b00110100110100000111: color_data = 12'b111011101110;
20'b00110100110100001000: color_data = 12'b111011101110;
20'b00110100110100001001: color_data = 12'b111111111111;
20'b00110100110100001010: color_data = 12'b111011101110;
20'b00110100110100001011: color_data = 12'b111011101110;
20'b00110100110100001101: color_data = 12'b111011101110;
20'b00110100110100001110: color_data = 12'b111011101110;
20'b00110100110100001111: color_data = 12'b111011101110;
20'b00110100110100010000: color_data = 12'b111011101110;
20'b00110100110100010111: color_data = 12'b111011101110;
20'b00110100110100011000: color_data = 12'b111011101110;
20'b00110100110100011001: color_data = 12'b111111111111;
20'b00110100110100011010: color_data = 12'b111111111111;
20'b00110100110100011011: color_data = 12'b111011101110;
20'b00110100110100011101: color_data = 12'b111011101110;
20'b00110100110100011110: color_data = 12'b111011101110;
20'b00110100110100011111: color_data = 12'b111011101110;
20'b00110100110100100000: color_data = 12'b111111111111;
20'b00110100110100100001: color_data = 12'b111011101110;
20'b00110100110100110011: color_data = 12'b111111111111;
20'b00110100110100110100: color_data = 12'b111011101110;
20'b00110100110100110101: color_data = 12'b111011101110;
20'b00110100110100110110: color_data = 12'b111011101110;
20'b00110100110100110111: color_data = 12'b111011101110;
20'b00110100110100111001: color_data = 12'b111011101110;
20'b00110100110100111010: color_data = 12'b111011101110;
20'b00110100110100111011: color_data = 12'b111011101110;
20'b00110100110100111100: color_data = 12'b111011101110;
20'b00110100110101000011: color_data = 12'b111011101110;
20'b00110100110101000100: color_data = 12'b111011101110;
20'b00110100110101000101: color_data = 12'b111011101110;
20'b00110100110101000110: color_data = 12'b111011101110;
20'b00110100110101000111: color_data = 12'b111011101110;
20'b00110100110101001001: color_data = 12'b111011101110;
20'b00110100110101001010: color_data = 12'b111011101110;
20'b00110100110101001011: color_data = 12'b111011101110;
20'b00110100110101001100: color_data = 12'b111111111111;
20'b00110100110101001101: color_data = 12'b111011101110;
20'b00110100110101011111: color_data = 12'b111011101110;
20'b00110100110101100000: color_data = 12'b111011101110;
20'b00110100110101100001: color_data = 12'b111011101110;
20'b00110100110101100010: color_data = 12'b111111111111;
20'b00110100110101100100: color_data = 12'b111011101110;
20'b00110100110101100101: color_data = 12'b111011101110;
20'b00110100110101100110: color_data = 12'b111011101110;
20'b00110100110101100111: color_data = 12'b111011101110;
20'b00110100110101101000: color_data = 12'b111011101110;
20'b00110100110101101111: color_data = 12'b111011101110;
20'b00110100110101110000: color_data = 12'b111011101110;
20'b00110100110101110001: color_data = 12'b111011101110;
20'b00110100110101110010: color_data = 12'b111011101110;
20'b00110100110101110011: color_data = 12'b111011101110;
20'b00110100110101110101: color_data = 12'b111111111111;
20'b00110100110101110110: color_data = 12'b111011101110;
20'b00110100110101110111: color_data = 12'b111011101110;
20'b00110100110101111000: color_data = 12'b111011101110;
20'b00110100110101111001: color_data = 12'b111011101110;
20'b00110101000100010111: color_data = 12'b111011101110;
20'b00110101000100011000: color_data = 12'b111011101110;
20'b00110101000100011001: color_data = 12'b111011101110;
20'b00110101000100011010: color_data = 12'b111011101110;
20'b00110101000100011011: color_data = 12'b111011101110;
20'b00110101000100011101: color_data = 12'b111011101110;
20'b00110101000100011110: color_data = 12'b111011101110;
20'b00110101000100011111: color_data = 12'b111011101110;
20'b00110101000100100000: color_data = 12'b111011101110;
20'b00110101000100100001: color_data = 12'b111111111111;
20'b00110101000100110011: color_data = 12'b111011101110;
20'b00110101000100110100: color_data = 12'b111011101110;
20'b00110101000100110101: color_data = 12'b111111111111;
20'b00110101000100110110: color_data = 12'b111011101110;
20'b00110101000100110111: color_data = 12'b111011101110;
20'b00110101000100111001: color_data = 12'b111011101110;
20'b00110101000100111010: color_data = 12'b111011101110;
20'b00110101000100111011: color_data = 12'b111011101110;
20'b00110101000100111100: color_data = 12'b111011101110;
20'b00110101000101000011: color_data = 12'b111011101110;
20'b00110101000101000100: color_data = 12'b111011101110;
20'b00110101000101000101: color_data = 12'b111011101110;
20'b00110101000101000110: color_data = 12'b111011101110;
20'b00110101000101000111: color_data = 12'b111011101110;
20'b00110101000101001001: color_data = 12'b111111111111;
20'b00110101000101001010: color_data = 12'b111011101110;
20'b00110101000101001011: color_data = 12'b111111111111;
20'b00110101000101001100: color_data = 12'b111011101110;
20'b00110101000101001101: color_data = 12'b111011101110;
20'b00110101000101011111: color_data = 12'b111011101110;
20'b00110101000101100000: color_data = 12'b111011101110;
20'b00110101000101100001: color_data = 12'b111011101110;
20'b00110101000101100010: color_data = 12'b111011101110;
20'b00110101000101100100: color_data = 12'b111011101110;
20'b00110101000101100101: color_data = 12'b111011101110;
20'b00110101000101100110: color_data = 12'b111011101110;
20'b00110101000101100111: color_data = 12'b111011101110;
20'b00110101000101101000: color_data = 12'b111011101110;
20'b00110101000101101111: color_data = 12'b111011101110;
20'b00110101000101110000: color_data = 12'b111011101110;
20'b00110101000101110001: color_data = 12'b111011101110;
20'b00110101000101110010: color_data = 12'b111011101110;
20'b00110101000101110011: color_data = 12'b111011101110;
20'b00110101000101110101: color_data = 12'b111011101110;
20'b00110101000101110110: color_data = 12'b111011101110;
20'b00110101000101110111: color_data = 12'b111011101110;
20'b00110101000101111000: color_data = 12'b111011101110;
20'b00110101000101111001: color_data = 12'b111011101110;
20'b00110101010011101011: color_data = 12'b111011101110;
20'b00110101010011101100: color_data = 12'b111011101110;
20'b00110101010011101101: color_data = 12'b111111111111;
20'b00110101010011101110: color_data = 12'b111011101110;
20'b00110101010011101111: color_data = 12'b111011101110;
20'b00110101010011110001: color_data = 12'b111111111111;
20'b00110101010011110010: color_data = 12'b111011101110;
20'b00110101010011110011: color_data = 12'b111011101110;
20'b00110101010011110100: color_data = 12'b111111111111;
20'b00110101010011110101: color_data = 12'b111011101110;
20'b00110101010011110111: color_data = 12'b111111111111;
20'b00110101010011111000: color_data = 12'b111111111111;
20'b00110101010011111001: color_data = 12'b111011101110;
20'b00110101010011111010: color_data = 12'b111011101110;
20'b00110101010011111100: color_data = 12'b111011101110;
20'b00110101010011111101: color_data = 12'b111011101110;
20'b00110101010011111110: color_data = 12'b111011101110;
20'b00110101010011111111: color_data = 12'b111011101110;
20'b00110101010100000001: color_data = 12'b111111111111;
20'b00110101010100000010: color_data = 12'b111011101110;
20'b00110101010100000011: color_data = 12'b111011101110;
20'b00110101010100000100: color_data = 12'b111011101110;
20'b00110101010100000101: color_data = 12'b111011101110;
20'b00110101010100000111: color_data = 12'b111011101110;
20'b00110101010100001000: color_data = 12'b111011101110;
20'b00110101010100001001: color_data = 12'b111111111111;
20'b00110101010100001010: color_data = 12'b111011101110;
20'b00110101010100001011: color_data = 12'b111011101110;
20'b00110101010100001101: color_data = 12'b111011101110;
20'b00110101010100001110: color_data = 12'b111011101110;
20'b00110101010100001111: color_data = 12'b111011101110;
20'b00110101010100010000: color_data = 12'b111011101110;
20'b00110101100011101011: color_data = 12'b111011101110;
20'b00110101100011101100: color_data = 12'b111011101110;
20'b00110101100011101101: color_data = 12'b111011101110;
20'b00110101100011101110: color_data = 12'b111111111111;
20'b00110101100011101111: color_data = 12'b111011101110;
20'b00110101100011110001: color_data = 12'b111011101110;
20'b00110101100011110010: color_data = 12'b111011101110;
20'b00110101100011110011: color_data = 12'b111111111111;
20'b00110101100011110100: color_data = 12'b111011101110;
20'b00110101100011110101: color_data = 12'b111011101110;
20'b00110101100011110111: color_data = 12'b111011101110;
20'b00110101100011111000: color_data = 12'b111011101110;
20'b00110101100011111001: color_data = 12'b111011101110;
20'b00110101100011111010: color_data = 12'b111011101110;
20'b00110101100011111100: color_data = 12'b111111111111;
20'b00110101100011111101: color_data = 12'b111111111111;
20'b00110101100011111110: color_data = 12'b111011101110;
20'b00110101100011111111: color_data = 12'b111011101110;
20'b00110101100100000001: color_data = 12'b111011101110;
20'b00110101100100000010: color_data = 12'b111011101110;
20'b00110101100100000011: color_data = 12'b111011101110;
20'b00110101100100000100: color_data = 12'b111011101110;
20'b00110101100100000101: color_data = 12'b111011101110;
20'b00110101100100000111: color_data = 12'b111011101110;
20'b00110101100100001000: color_data = 12'b111011101110;
20'b00110101100100001001: color_data = 12'b111011101110;
20'b00110101100100001010: color_data = 12'b111111111111;
20'b00110101100100001011: color_data = 12'b111011101110;
20'b00110101100100001101: color_data = 12'b111111111111;
20'b00110101100100001110: color_data = 12'b111011101110;
20'b00110101100100001111: color_data = 12'b111011101110;
20'b00110101100100010000: color_data = 12'b111011101110;
20'b00110101100100010111: color_data = 12'b111011101110;
20'b00110101100100011000: color_data = 12'b111011101110;
20'b00110101100100011001: color_data = 12'b111011101110;
20'b00110101100100011010: color_data = 12'b111011101110;
20'b00110101100100011011: color_data = 12'b111011101110;
20'b00110101100100011101: color_data = 12'b111111111111;
20'b00110101100100011110: color_data = 12'b111011101110;
20'b00110101100100011111: color_data = 12'b111111111111;
20'b00110101100100100000: color_data = 12'b111011101110;
20'b00110101100100100001: color_data = 12'b111011101110;
20'b00110101100100110011: color_data = 12'b111011101110;
20'b00110101100100110100: color_data = 12'b111011101110;
20'b00110101100100110101: color_data = 12'b111011101110;
20'b00110101100100110110: color_data = 12'b111111111111;
20'b00110101100100110111: color_data = 12'b111011101110;
20'b00110101100100111001: color_data = 12'b111011101110;
20'b00110101100100111010: color_data = 12'b111011101110;
20'b00110101100100111011: color_data = 12'b111011101110;
20'b00110101100100111100: color_data = 12'b111111111111;
20'b00110101100101000011: color_data = 12'b111011101110;
20'b00110101100101000100: color_data = 12'b111011101110;
20'b00110101100101000101: color_data = 12'b111011101110;
20'b00110101100101000110: color_data = 12'b111011101110;
20'b00110101100101000111: color_data = 12'b111011101110;
20'b00110101100101001001: color_data = 12'b111111111111;
20'b00110101100101001010: color_data = 12'b111011101110;
20'b00110101100101001011: color_data = 12'b111011101110;
20'b00110101100101001100: color_data = 12'b111011101110;
20'b00110101100101001101: color_data = 12'b111011101110;
20'b00110101100101011111: color_data = 12'b111011101110;
20'b00110101100101100000: color_data = 12'b111011101110;
20'b00110101100101100001: color_data = 12'b111011101110;
20'b00110101100101100010: color_data = 12'b111011101110;
20'b00110101100101100100: color_data = 12'b111011101110;
20'b00110101100101100101: color_data = 12'b111011101110;
20'b00110101100101100110: color_data = 12'b111011101110;
20'b00110101100101100111: color_data = 12'b111011101110;
20'b00110101100101101000: color_data = 12'b111011101110;
20'b00110101100101101111: color_data = 12'b111011101110;
20'b00110101100101110000: color_data = 12'b111011101110;
20'b00110101100101110001: color_data = 12'b111011101110;
20'b00110101100101110010: color_data = 12'b111011101110;
20'b00110101100101110011: color_data = 12'b111011101110;
20'b00110101100101110101: color_data = 12'b111011101110;
20'b00110101100101110110: color_data = 12'b111011101110;
20'b00110101100101110111: color_data = 12'b111011101110;
20'b00110101100101111000: color_data = 12'b111011101110;
20'b00110101100101111001: color_data = 12'b111011101110;
20'b00110101100101111011: color_data = 12'b111011101110;
20'b00110101100101111100: color_data = 12'b111011101110;
20'b00110101100101111101: color_data = 12'b111011101110;
20'b00110101100101111110: color_data = 12'b111011101110;
20'b00110101100110000000: color_data = 12'b111011101110;
20'b00110101100110000001: color_data = 12'b111111111111;
20'b00110101100110000010: color_data = 12'b111011101110;
20'b00110101100110000011: color_data = 12'b111011101110;
20'b00110101100110000100: color_data = 12'b111011101110;
20'b00110101100110000110: color_data = 12'b111011101110;
20'b00110101100110000111: color_data = 12'b111011101110;
20'b00110101100110001000: color_data = 12'b111011101110;
20'b00110101100110001001: color_data = 12'b111011101110;
20'b00110101100110001011: color_data = 12'b111011101110;
20'b00110101100110001100: color_data = 12'b111011101110;
20'b00110101100110001101: color_data = 12'b111011101110;
20'b00110101100110001110: color_data = 12'b111111111111;
20'b00110101100110001111: color_data = 12'b111011101110;
20'b00110101100110010001: color_data = 12'b111011101110;
20'b00110101100110010010: color_data = 12'b111011101110;
20'b00110101100110010011: color_data = 12'b111111111111;
20'b00110101100110010100: color_data = 12'b111011101110;
20'b00110101110011101011: color_data = 12'b111011101110;
20'b00110101110011101100: color_data = 12'b111011101110;
20'b00110101110011101101: color_data = 12'b111011101110;
20'b00110101110011101110: color_data = 12'b111011101110;
20'b00110101110011101111: color_data = 12'b111011101110;
20'b00110101110011110001: color_data = 12'b111011101110;
20'b00110101110011110010: color_data = 12'b111111111111;
20'b00110101110011110011: color_data = 12'b111011101110;
20'b00110101110011110100: color_data = 12'b111011101110;
20'b00110101110011110101: color_data = 12'b111011101110;
20'b00110101110011110111: color_data = 12'b111011101110;
20'b00110101110011111000: color_data = 12'b111011101110;
20'b00110101110011111001: color_data = 12'b111011101110;
20'b00110101110011111010: color_data = 12'b111011101110;
20'b00110101110011111100: color_data = 12'b111011101110;
20'b00110101110011111101: color_data = 12'b111011101110;
20'b00110101110011111110: color_data = 12'b111011101110;
20'b00110101110011111111: color_data = 12'b111011101110;
20'b00110101110100000001: color_data = 12'b111011101110;
20'b00110101110100000010: color_data = 12'b111111111111;
20'b00110101110100000011: color_data = 12'b111011101110;
20'b00110101110100000100: color_data = 12'b111011101110;
20'b00110101110100000101: color_data = 12'b111111111111;
20'b00110101110100000111: color_data = 12'b111011101110;
20'b00110101110100001000: color_data = 12'b111011101110;
20'b00110101110100001001: color_data = 12'b111011101110;
20'b00110101110100001010: color_data = 12'b111011101110;
20'b00110101110100001011: color_data = 12'b111011101110;
20'b00110101110100001101: color_data = 12'b111011101110;
20'b00110101110100001110: color_data = 12'b111011101110;
20'b00110101110100001111: color_data = 12'b111111111111;
20'b00110101110100010000: color_data = 12'b111011101110;
20'b00110101110100010111: color_data = 12'b111011101110;
20'b00110101110100011000: color_data = 12'b111011101110;
20'b00110101110100011001: color_data = 12'b111011101110;
20'b00110101110100011010: color_data = 12'b111011101110;
20'b00110101110100011011: color_data = 12'b111011101110;
20'b00110101110100011101: color_data = 12'b111011101110;
20'b00110101110100011110: color_data = 12'b111011101110;
20'b00110101110100011111: color_data = 12'b111011101110;
20'b00110101110100100000: color_data = 12'b111011101110;
20'b00110101110100100001: color_data = 12'b111011101110;
20'b00110101110100110011: color_data = 12'b111011101110;
20'b00110101110100110100: color_data = 12'b111011101110;
20'b00110101110100110101: color_data = 12'b111011101110;
20'b00110101110100110110: color_data = 12'b111011101110;
20'b00110101110100110111: color_data = 12'b111011101110;
20'b00110101110100111001: color_data = 12'b111011101110;
20'b00110101110100111010: color_data = 12'b111011101110;
20'b00110101110100111011: color_data = 12'b111011101110;
20'b00110101110100111100: color_data = 12'b111011101110;
20'b00110101110101000011: color_data = 12'b111011101110;
20'b00110101110101000100: color_data = 12'b111011101110;
20'b00110101110101000101: color_data = 12'b111011101110;
20'b00110101110101000110: color_data = 12'b111011101110;
20'b00110101110101000111: color_data = 12'b111011101110;
20'b00110101110101001001: color_data = 12'b111011101110;
20'b00110101110101001010: color_data = 12'b111011101110;
20'b00110101110101001011: color_data = 12'b111011101110;
20'b00110101110101001100: color_data = 12'b111011101110;
20'b00110101110101001101: color_data = 12'b111011101110;
20'b00110101110101011111: color_data = 12'b111011101110;
20'b00110101110101100000: color_data = 12'b111011101110;
20'b00110101110101100001: color_data = 12'b111011101110;
20'b00110101110101100010: color_data = 12'b111011101110;
20'b00110101110101100100: color_data = 12'b111011101110;
20'b00110101110101100101: color_data = 12'b111111111111;
20'b00110101110101100110: color_data = 12'b111011101110;
20'b00110101110101100111: color_data = 12'b111011101110;
20'b00110101110101101000: color_data = 12'b111011101110;
20'b00110101110101101111: color_data = 12'b111011101110;
20'b00110101110101110000: color_data = 12'b111011101110;
20'b00110101110101110001: color_data = 12'b111011101110;
20'b00110101110101110010: color_data = 12'b111111111111;
20'b00110101110101110011: color_data = 12'b111011101110;
20'b00110101110101110101: color_data = 12'b111011101110;
20'b00110101110101110110: color_data = 12'b111011101110;
20'b00110101110101110111: color_data = 12'b111011101110;
20'b00110101110101111000: color_data = 12'b111011101110;
20'b00110101110101111001: color_data = 12'b111011101110;
20'b00110101110101111011: color_data = 12'b111011101110;
20'b00110101110101111100: color_data = 12'b111011101110;
20'b00110101110101111101: color_data = 12'b111011101110;
20'b00110101110101111110: color_data = 12'b111011101110;
20'b00110101110110000000: color_data = 12'b111011101110;
20'b00110101110110000001: color_data = 12'b111011101110;
20'b00110101110110000010: color_data = 12'b111011101110;
20'b00110101110110000011: color_data = 12'b111011101110;
20'b00110101110110000100: color_data = 12'b111011101110;
20'b00110101110110000110: color_data = 12'b111011101110;
20'b00110101110110000111: color_data = 12'b111011101110;
20'b00110101110110001000: color_data = 12'b111011101110;
20'b00110101110110001001: color_data = 12'b111011101110;
20'b00110101110110001011: color_data = 12'b111011101110;
20'b00110101110110001100: color_data = 12'b111011101110;
20'b00110101110110001101: color_data = 12'b111011101110;
20'b00110101110110001110: color_data = 12'b111011101110;
20'b00110101110110001111: color_data = 12'b111011101110;
20'b00110101110110010001: color_data = 12'b111011101110;
20'b00110101110110010010: color_data = 12'b111011101110;
20'b00110101110110010011: color_data = 12'b111011101110;
20'b00110101110110010100: color_data = 12'b111011101110;
20'b00110110000011101011: color_data = 12'b111011101110;
20'b00110110000011101100: color_data = 12'b111011101110;
20'b00110110000011101101: color_data = 12'b111011101110;
20'b00110110000011101110: color_data = 12'b111011101110;
20'b00110110000011101111: color_data = 12'b111011101110;
20'b00110110000011110001: color_data = 12'b111011101110;
20'b00110110000011110010: color_data = 12'b111011101110;
20'b00110110000011110011: color_data = 12'b111011101110;
20'b00110110000011110100: color_data = 12'b111011101110;
20'b00110110000011110101: color_data = 12'b111011101110;
20'b00110110000011110111: color_data = 12'b111011101110;
20'b00110110000011111000: color_data = 12'b111011101110;
20'b00110110000011111001: color_data = 12'b111011101110;
20'b00110110000011111010: color_data = 12'b111011101110;
20'b00110110000011111100: color_data = 12'b111011101110;
20'b00110110000011111101: color_data = 12'b111111111111;
20'b00110110000011111110: color_data = 12'b111011101110;
20'b00110110000011111111: color_data = 12'b111011101110;
20'b00110110000100000001: color_data = 12'b111011101110;
20'b00110110000100000010: color_data = 12'b111011101110;
20'b00110110000100000011: color_data = 12'b111011101110;
20'b00110110000100000100: color_data = 12'b111011101110;
20'b00110110000100000101: color_data = 12'b111011101110;
20'b00110110000100000111: color_data = 12'b111011101110;
20'b00110110000100001000: color_data = 12'b111011101110;
20'b00110110000100001001: color_data = 12'b111111111111;
20'b00110110000100001010: color_data = 12'b111011101110;
20'b00110110000100001011: color_data = 12'b111011101110;
20'b00110110000100001101: color_data = 12'b111011101110;
20'b00110110000100001110: color_data = 12'b111011101110;
20'b00110110000100001111: color_data = 12'b111011101110;
20'b00110110000100010000: color_data = 12'b111011101110;
20'b00110110000100010111: color_data = 12'b111011101110;
20'b00110110000100011000: color_data = 12'b111011101110;
20'b00110110000100011001: color_data = 12'b111011101110;
20'b00110110000100011010: color_data = 12'b111111111111;
20'b00110110000100011011: color_data = 12'b111011101110;
20'b00110110000100011101: color_data = 12'b111011101110;
20'b00110110000100011110: color_data = 12'b111011101110;
20'b00110110000100011111: color_data = 12'b111011101110;
20'b00110110000100100000: color_data = 12'b111011101110;
20'b00110110000100100001: color_data = 12'b111011101110;
20'b00110110000100110011: color_data = 12'b111011101110;
20'b00110110000100110100: color_data = 12'b111011101110;
20'b00110110000100110101: color_data = 12'b111011101110;
20'b00110110000100110110: color_data = 12'b111011101110;
20'b00110110000100110111: color_data = 12'b111011101110;
20'b00110110000100111001: color_data = 12'b111011101110;
20'b00110110000100111010: color_data = 12'b111011101110;
20'b00110110000100111011: color_data = 12'b111011101110;
20'b00110110000100111100: color_data = 12'b111011101110;
20'b00110110000101000011: color_data = 12'b111011101110;
20'b00110110000101000100: color_data = 12'b111011101110;
20'b00110110000101000101: color_data = 12'b111011101110;
20'b00110110000101000110: color_data = 12'b111011101110;
20'b00110110000101000111: color_data = 12'b111011101110;
20'b00110110000101001001: color_data = 12'b111011101110;
20'b00110110000101001010: color_data = 12'b111011101110;
20'b00110110000101001011: color_data = 12'b111011101110;
20'b00110110000101001100: color_data = 12'b111011101110;
20'b00110110000101001101: color_data = 12'b111011101110;
20'b00110110000101011111: color_data = 12'b111011101110;
20'b00110110000101100000: color_data = 12'b111011101110;
20'b00110110000101100001: color_data = 12'b111011101110;
20'b00110110000101100010: color_data = 12'b111011101110;
20'b00110110000101100100: color_data = 12'b111011101110;
20'b00110110000101100101: color_data = 12'b111111111111;
20'b00110110000101100110: color_data = 12'b111011101110;
20'b00110110000101100111: color_data = 12'b111011101110;
20'b00110110000101101000: color_data = 12'b111011101110;
20'b00110110000101101111: color_data = 12'b111011101110;
20'b00110110000101110000: color_data = 12'b111011101110;
20'b00110110000101110001: color_data = 12'b111011101110;
20'b00110110000101110010: color_data = 12'b111111111111;
20'b00110110000101110011: color_data = 12'b111011101110;
20'b00110110000101110101: color_data = 12'b111011101110;
20'b00110110000101110110: color_data = 12'b111011101110;
20'b00110110000101110111: color_data = 12'b111011101110;
20'b00110110000101111000: color_data = 12'b111011101110;
20'b00110110000101111001: color_data = 12'b111011101110;
20'b00110110000101111011: color_data = 12'b111111111111;
20'b00110110000101111100: color_data = 12'b111011101110;
20'b00110110000101111101: color_data = 12'b111011101110;
20'b00110110000101111110: color_data = 12'b111011101110;
20'b00110110000110000000: color_data = 12'b111011101110;
20'b00110110000110000001: color_data = 12'b111011101110;
20'b00110110000110000010: color_data = 12'b111011101110;
20'b00110110000110000011: color_data = 12'b111011101110;
20'b00110110000110000100: color_data = 12'b111011101110;
20'b00110110000110000110: color_data = 12'b111011101110;
20'b00110110000110000111: color_data = 12'b111111111111;
20'b00110110000110001000: color_data = 12'b111111111111;
20'b00110110000110001001: color_data = 12'b111011101110;
20'b00110110000110001011: color_data = 12'b111011101110;
20'b00110110000110001100: color_data = 12'b111011101110;
20'b00110110000110001101: color_data = 12'b111011101110;
20'b00110110000110001110: color_data = 12'b111011101110;
20'b00110110000110001111: color_data = 12'b111011101110;
20'b00110110000110010001: color_data = 12'b111011101110;
20'b00110110000110010010: color_data = 12'b111011101110;
20'b00110110000110010011: color_data = 12'b111011101110;
20'b00110110000110010100: color_data = 12'b111011101110;
20'b00110110010011101011: color_data = 12'b111011101110;
20'b00110110010011101100: color_data = 12'b111011101110;
20'b00110110010011101101: color_data = 12'b111011101110;
20'b00110110010011101110: color_data = 12'b111011101110;
20'b00110110010011101111: color_data = 12'b111011101110;
20'b00110110010011110001: color_data = 12'b111011101110;
20'b00110110010011110010: color_data = 12'b111011101110;
20'b00110110010011110011: color_data = 12'b111011101110;
20'b00110110010011110100: color_data = 12'b111011101110;
20'b00110110010011110101: color_data = 12'b111011101110;
20'b00110110010011110111: color_data = 12'b111011101110;
20'b00110110010011111000: color_data = 12'b111011101110;
20'b00110110010011111001: color_data = 12'b111011101110;
20'b00110110010011111010: color_data = 12'b111011101110;
20'b00110110010011111100: color_data = 12'b111011101110;
20'b00110110010011111101: color_data = 12'b111011101110;
20'b00110110010011111110: color_data = 12'b111011101110;
20'b00110110010011111111: color_data = 12'b111011101110;
20'b00110110010100000001: color_data = 12'b111011101110;
20'b00110110010100000010: color_data = 12'b111011101110;
20'b00110110010100000011: color_data = 12'b111011101110;
20'b00110110010100000100: color_data = 12'b111011101110;
20'b00110110010100000101: color_data = 12'b111011101110;
20'b00110110010100000111: color_data = 12'b111011101110;
20'b00110110010100001000: color_data = 12'b111011101110;
20'b00110110010100001001: color_data = 12'b111011101110;
20'b00110110010100001010: color_data = 12'b111011101110;
20'b00110110010100001011: color_data = 12'b111011101110;
20'b00110110010100001101: color_data = 12'b111111111111;
20'b00110110010100001110: color_data = 12'b111011101110;
20'b00110110010100001111: color_data = 12'b111011101110;
20'b00110110010100010000: color_data = 12'b111011101110;
20'b00110110010100010111: color_data = 12'b111011101110;
20'b00110110010100011000: color_data = 12'b111011101110;
20'b00110110010100011001: color_data = 12'b111011101110;
20'b00110110010100011010: color_data = 12'b111011101110;
20'b00110110010100011011: color_data = 12'b111011101110;
20'b00110110010100011101: color_data = 12'b111011101110;
20'b00110110010100011110: color_data = 12'b111011101110;
20'b00110110010100011111: color_data = 12'b111011101110;
20'b00110110010100100000: color_data = 12'b111011101110;
20'b00110110010100100001: color_data = 12'b111011101110;
20'b00110110010100110011: color_data = 12'b111011101110;
20'b00110110010100110100: color_data = 12'b111011101110;
20'b00110110010100110101: color_data = 12'b111011101110;
20'b00110110010100110110: color_data = 12'b111011101110;
20'b00110110010100110111: color_data = 12'b111011101110;
20'b00110110010100111001: color_data = 12'b111011101110;
20'b00110110010100111010: color_data = 12'b111111111111;
20'b00110110010100111011: color_data = 12'b111011101110;
20'b00110110010100111100: color_data = 12'b111011101110;
20'b00110110010101000011: color_data = 12'b111011101110;
20'b00110110010101000100: color_data = 12'b111011101110;
20'b00110110010101000101: color_data = 12'b111011101110;
20'b00110110010101000110: color_data = 12'b111011101110;
20'b00110110010101000111: color_data = 12'b111011101110;
20'b00110110010101001001: color_data = 12'b111111111111;
20'b00110110010101001010: color_data = 12'b111011101110;
20'b00110110010101001011: color_data = 12'b111011101110;
20'b00110110010101001100: color_data = 12'b111011101110;
20'b00110110010101001101: color_data = 12'b111011101110;
20'b00110110010101011111: color_data = 12'b111011101110;
20'b00110110010101100000: color_data = 12'b111011101110;
20'b00110110010101100001: color_data = 12'b111011101110;
20'b00110110010101100010: color_data = 12'b111011101110;
20'b00110110010101100100: color_data = 12'b111011101110;
20'b00110110010101100101: color_data = 12'b111011101110;
20'b00110110010101100110: color_data = 12'b111011101110;
20'b00110110010101100111: color_data = 12'b111011101110;
20'b00110110010101101000: color_data = 12'b111011101110;
20'b00110110010101101111: color_data = 12'b111011101110;
20'b00110110010101110000: color_data = 12'b111011101110;
20'b00110110010101110001: color_data = 12'b111011101110;
20'b00110110010101110010: color_data = 12'b111011101110;
20'b00110110010101110011: color_data = 12'b111011101110;
20'b00110110010101110101: color_data = 12'b111011101110;
20'b00110110010101110110: color_data = 12'b111011101110;
20'b00110110010101110111: color_data = 12'b111011101110;
20'b00110110010101111000: color_data = 12'b111011101110;
20'b00110110010101111001: color_data = 12'b111011101110;
20'b00110110010101111011: color_data = 12'b111011101110;
20'b00110110010101111100: color_data = 12'b111011101110;
20'b00110110010101111101: color_data = 12'b111011101110;
20'b00110110010101111110: color_data = 12'b111111111111;
20'b00110110010110000000: color_data = 12'b111011101110;
20'b00110110010110000001: color_data = 12'b111011101110;
20'b00110110010110000010: color_data = 12'b111011101110;
20'b00110110010110000011: color_data = 12'b111011101110;
20'b00110110010110000100: color_data = 12'b111011101110;
20'b00110110010110000110: color_data = 12'b111111111111;
20'b00110110010110000111: color_data = 12'b111011101110;
20'b00110110010110001000: color_data = 12'b111011101110;
20'b00110110010110001001: color_data = 12'b111111111111;
20'b00110110010110001011: color_data = 12'b111011101110;
20'b00110110010110001100: color_data = 12'b111011101110;
20'b00110110010110001101: color_data = 12'b111011101110;
20'b00110110010110001110: color_data = 12'b111011101110;
20'b00110110010110001111: color_data = 12'b111011101110;
20'b00110110010110010001: color_data = 12'b111011101110;
20'b00110110010110010010: color_data = 12'b111111111111;
20'b00110110010110010011: color_data = 12'b111011101110;
20'b00110110010110010100: color_data = 12'b111011101110;
20'b00110110110011110001: color_data = 12'b111011101110;
20'b00110110110011110010: color_data = 12'b111011101110;
20'b00110110110011110011: color_data = 12'b111011101110;
20'b00110110110011110100: color_data = 12'b111011101110;
20'b00110110110011110101: color_data = 12'b111011101110;
20'b00110110110011110111: color_data = 12'b111011101110;
20'b00110110110011111000: color_data = 12'b111011101110;
20'b00110110110011111001: color_data = 12'b111011101110;
20'b00110110110011111010: color_data = 12'b111011101110;
20'b00110110110011111100: color_data = 12'b111011101110;
20'b00110110110011111101: color_data = 12'b111011101110;
20'b00110110110011111110: color_data = 12'b111011101110;
20'b00110110110011111111: color_data = 12'b111011101110;
20'b00110110110100000001: color_data = 12'b111011101110;
20'b00110110110100000010: color_data = 12'b111011101110;
20'b00110110110100000011: color_data = 12'b111011101110;
20'b00110110110100000100: color_data = 12'b111011101110;
20'b00110110110100000101: color_data = 12'b111011101110;
20'b00110110110100000111: color_data = 12'b111011101110;
20'b00110110110100001000: color_data = 12'b111011101110;
20'b00110110110100001001: color_data = 12'b111011101110;
20'b00110110110100001010: color_data = 12'b111011101110;
20'b00110110110100001011: color_data = 12'b111011101110;
20'b00110110110100010111: color_data = 12'b111011101110;
20'b00110110110100011000: color_data = 12'b111011101110;
20'b00110110110100011001: color_data = 12'b111011101110;
20'b00110110110100011010: color_data = 12'b111011101110;
20'b00110110110100011011: color_data = 12'b111011101110;
20'b00110110110100011101: color_data = 12'b111011101110;
20'b00110110110100011110: color_data = 12'b111011101110;
20'b00110110110100011111: color_data = 12'b111011101110;
20'b00110110110100100000: color_data = 12'b111011101110;
20'b00110110110100100001: color_data = 12'b111111111111;
20'b00110110110100110011: color_data = 12'b111011101110;
20'b00110110110100110100: color_data = 12'b111011101110;
20'b00110110110100110101: color_data = 12'b111011101110;
20'b00110110110100110110: color_data = 12'b111011101110;
20'b00110110110100110111: color_data = 12'b111011101110;
20'b00110110110100111001: color_data = 12'b111011101110;
20'b00110110110100111010: color_data = 12'b111111111111;
20'b00110110110100111011: color_data = 12'b111111111111;
20'b00110110110100111100: color_data = 12'b111011101110;
20'b00110110110101000011: color_data = 12'b111011101110;
20'b00110110110101000100: color_data = 12'b111011101110;
20'b00110110110101000101: color_data = 12'b111011101110;
20'b00110110110101000110: color_data = 12'b111011101110;
20'b00110110110101000111: color_data = 12'b111011101110;
20'b00110110110101001001: color_data = 12'b111111111111;
20'b00110110110101001010: color_data = 12'b111011101110;
20'b00110110110101001011: color_data = 12'b111111111111;
20'b00110110110101001100: color_data = 12'b111011101110;
20'b00110110110101001101: color_data = 12'b111011101110;
20'b00110110110101011111: color_data = 12'b111011101110;
20'b00110110110101100000: color_data = 12'b111011101110;
20'b00110110110101100001: color_data = 12'b111011101110;
20'b00110110110101100010: color_data = 12'b111011101110;
20'b00110110110101100100: color_data = 12'b111011101110;
20'b00110110110101100101: color_data = 12'b111011101110;
20'b00110110110101100110: color_data = 12'b111011101110;
20'b00110110110101100111: color_data = 12'b111011101110;
20'b00110110110101101000: color_data = 12'b111011101110;
20'b00110110110101101111: color_data = 12'b111011101110;
20'b00110110110101110000: color_data = 12'b111011101110;
20'b00110110110101110001: color_data = 12'b111011101110;
20'b00110110110101110010: color_data = 12'b111011101110;
20'b00110110110101110011: color_data = 12'b111011101110;
20'b00110110110101110101: color_data = 12'b111011101110;
20'b00110110110101110110: color_data = 12'b111011101110;
20'b00110110110101110111: color_data = 12'b111011101110;
20'b00110110110101111000: color_data = 12'b111011101110;
20'b00110110110101111001: color_data = 12'b111011101110;
20'b00110110110101111011: color_data = 12'b111011101110;
20'b00110110110101111100: color_data = 12'b111011101110;
20'b00110110110101111101: color_data = 12'b111111111111;
20'b00110110110101111110: color_data = 12'b111011101110;
20'b00110110110110000000: color_data = 12'b111011101110;
20'b00110110110110000001: color_data = 12'b111011101110;
20'b00110110110110000010: color_data = 12'b111111111111;
20'b00110110110110000011: color_data = 12'b111011101110;
20'b00110110110110000100: color_data = 12'b111011101110;
20'b00110110110110000110: color_data = 12'b111011101110;
20'b00110110110110000111: color_data = 12'b111011101110;
20'b00110110110110001000: color_data = 12'b111011101110;
20'b00110110110110001001: color_data = 12'b111011101110;
20'b00110110110110001011: color_data = 12'b111011101110;
20'b00110110110110001100: color_data = 12'b111011101110;
20'b00110110110110001101: color_data = 12'b111111111111;
20'b00110110110110001110: color_data = 12'b111011101110;
20'b00110110110110001111: color_data = 12'b111011101110;
20'b00110110110110010001: color_data = 12'b111011101110;
20'b00110110110110010010: color_data = 12'b111111111111;
20'b00110110110110010011: color_data = 12'b111111111111;
20'b00110110110110010100: color_data = 12'b111011101110;
20'b00110111000011110001: color_data = 12'b111011101110;
20'b00110111000011110010: color_data = 12'b111011101110;
20'b00110111000011110011: color_data = 12'b111111111111;
20'b00110111000011110100: color_data = 12'b111011101110;
20'b00110111000011110101: color_data = 12'b111011101110;
20'b00110111000011110111: color_data = 12'b111011101110;
20'b00110111000011111000: color_data = 12'b111011101110;
20'b00110111000011111001: color_data = 12'b111011101110;
20'b00110111000011111010: color_data = 12'b111111111111;
20'b00110111000011111100: color_data = 12'b111011101110;
20'b00110111000011111101: color_data = 12'b111011101110;
20'b00110111000011111110: color_data = 12'b111011101110;
20'b00110111000011111111: color_data = 12'b111011101110;
20'b00110111000100000001: color_data = 12'b111011101110;
20'b00110111000100000010: color_data = 12'b111011101110;
20'b00110111000100000011: color_data = 12'b111111111111;
20'b00110111000100000100: color_data = 12'b111011101110;
20'b00110111000100000101: color_data = 12'b111011101110;
20'b00110111000100000111: color_data = 12'b111011101110;
20'b00110111000100001000: color_data = 12'b111011101110;
20'b00110111000100001001: color_data = 12'b111011101110;
20'b00110111000100001010: color_data = 12'b111011101110;
20'b00110111000100001011: color_data = 12'b111111111111;
20'b00110111000100010111: color_data = 12'b111011101110;
20'b00110111000100011000: color_data = 12'b111011101110;
20'b00110111000100011001: color_data = 12'b111011101110;
20'b00110111000100011010: color_data = 12'b111011101110;
20'b00110111000100011011: color_data = 12'b111011101110;
20'b00110111000100011101: color_data = 12'b111111111111;
20'b00110111000100011110: color_data = 12'b111011101110;
20'b00110111000100011111: color_data = 12'b111011101110;
20'b00110111000100100000: color_data = 12'b111011101110;
20'b00110111000100100001: color_data = 12'b111011101110;
20'b00110111000100110011: color_data = 12'b111011101110;
20'b00110111000100110100: color_data = 12'b111011101110;
20'b00110111000100110101: color_data = 12'b111011101110;
20'b00110111000100110110: color_data = 12'b111011101110;
20'b00110111000100110111: color_data = 12'b111011101110;
20'b00110111000100111001: color_data = 12'b111011101110;
20'b00110111000100111010: color_data = 12'b111011101110;
20'b00110111000100111011: color_data = 12'b111011101110;
20'b00110111000100111100: color_data = 12'b111011101110;
20'b00110111000101000011: color_data = 12'b111011101110;
20'b00110111000101000100: color_data = 12'b111011101110;
20'b00110111000101000101: color_data = 12'b111011101110;
20'b00110111000101000110: color_data = 12'b111011101110;
20'b00110111000101000111: color_data = 12'b111011101110;
20'b00110111000101001001: color_data = 12'b111011101110;
20'b00110111000101001010: color_data = 12'b111011101110;
20'b00110111000101001011: color_data = 12'b111011101110;
20'b00110111000101001100: color_data = 12'b111111111111;
20'b00110111000101001101: color_data = 12'b111011101110;
20'b00110111000101011111: color_data = 12'b111011101110;
20'b00110111000101100000: color_data = 12'b111011101110;
20'b00110111000101100001: color_data = 12'b111011101110;
20'b00110111000101100010: color_data = 12'b111111111111;
20'b00110111000101100100: color_data = 12'b111011101110;
20'b00110111000101100101: color_data = 12'b111011101110;
20'b00110111000101100110: color_data = 12'b111011101110;
20'b00110111000101100111: color_data = 12'b111011101110;
20'b00110111000101101000: color_data = 12'b111011101110;
20'b00110111000101101111: color_data = 12'b111011101110;
20'b00110111000101110000: color_data = 12'b111011101110;
20'b00110111000101110001: color_data = 12'b111011101110;
20'b00110111000101110010: color_data = 12'b111011101110;
20'b00110111000101110011: color_data = 12'b111011101110;
20'b00110111000101110101: color_data = 12'b111111111111;
20'b00110111000101110110: color_data = 12'b111011101110;
20'b00110111000101110111: color_data = 12'b111011101110;
20'b00110111000101111000: color_data = 12'b111011101110;
20'b00110111000101111001: color_data = 12'b111011101110;
20'b00110111000101111011: color_data = 12'b111011101110;
20'b00110111000101111100: color_data = 12'b111011101110;
20'b00110111000101111101: color_data = 12'b111011101110;
20'b00110111000101111110: color_data = 12'b111011101110;
20'b00110111000110000000: color_data = 12'b111011101110;
20'b00110111000110000001: color_data = 12'b111011101110;
20'b00110111000110000010: color_data = 12'b111011101110;
20'b00110111000110000011: color_data = 12'b111011101110;
20'b00110111000110000100: color_data = 12'b111011101110;
20'b00110111000110000110: color_data = 12'b111011101110;
20'b00110111000110000111: color_data = 12'b111011101110;
20'b00110111000110001000: color_data = 12'b111011101110;
20'b00110111000110001001: color_data = 12'b111011101110;
20'b00110111000110001011: color_data = 12'b111011101110;
20'b00110111000110001100: color_data = 12'b111011101110;
20'b00110111000110001101: color_data = 12'b111011101110;
20'b00110111000110001110: color_data = 12'b111011101110;
20'b00110111000110001111: color_data = 12'b111011101110;
20'b00110111000110010001: color_data = 12'b111011101110;
20'b00110111000110010010: color_data = 12'b111011101110;
20'b00110111000110010011: color_data = 12'b111011101110;
20'b00110111000110010100: color_data = 12'b111011101110;
20'b00110111010011110001: color_data = 12'b111011101110;
20'b00110111010011110010: color_data = 12'b111011101110;
20'b00110111010011110011: color_data = 12'b111011101110;
20'b00110111010011110100: color_data = 12'b111111111111;
20'b00110111010011110101: color_data = 12'b111011101110;
20'b00110111010011110111: color_data = 12'b111011101110;
20'b00110111010011111000: color_data = 12'b111011101110;
20'b00110111010011111001: color_data = 12'b111011101110;
20'b00110111010011111010: color_data = 12'b111011101110;
20'b00110111010011111100: color_data = 12'b111111111111;
20'b00110111010011111101: color_data = 12'b111011101110;
20'b00110111010011111110: color_data = 12'b111011101110;
20'b00110111010011111111: color_data = 12'b111011101110;
20'b00110111010100000001: color_data = 12'b111011101110;
20'b00110111010100000010: color_data = 12'b111011101110;
20'b00110111010100000011: color_data = 12'b111011101110;
20'b00110111010100000100: color_data = 12'b111111111111;
20'b00110111010100000101: color_data = 12'b111011101110;
20'b00110111010100000111: color_data = 12'b111011101110;
20'b00110111010100001000: color_data = 12'b111011101110;
20'b00110111010100001001: color_data = 12'b111011101110;
20'b00110111010100001010: color_data = 12'b111011101110;
20'b00110111010100001011: color_data = 12'b111011101110;
20'b00110111010100010111: color_data = 12'b111011101110;
20'b00110111010100011000: color_data = 12'b111011101110;
20'b00110111010100011001: color_data = 12'b111011101110;
20'b00110111010100011010: color_data = 12'b111011101110;
20'b00110111010100011011: color_data = 12'b111111111111;
20'b00110111010100011101: color_data = 12'b111011101110;
20'b00110111010100011110: color_data = 12'b111011101110;
20'b00110111010100011111: color_data = 12'b111011101110;
20'b00110111010100100000: color_data = 12'b111011101110;
20'b00110111010100100001: color_data = 12'b111011101110;
20'b00110111010100110011: color_data = 12'b111011101110;
20'b00110111010100110100: color_data = 12'b111111111111;
20'b00110111010100110101: color_data = 12'b111011101110;
20'b00110111010100110110: color_data = 12'b111011101110;
20'b00110111010100110111: color_data = 12'b111011101110;
20'b00110111010100111001: color_data = 12'b111011101110;
20'b00110111010100111010: color_data = 12'b111111111111;
20'b00110111010100111011: color_data = 12'b111011101110;
20'b00110111010100111100: color_data = 12'b111011101110;
20'b00110111010101000011: color_data = 12'b111011101110;
20'b00110111010101000100: color_data = 12'b111111111111;
20'b00110111010101000101: color_data = 12'b111011101110;
20'b00110111010101000110: color_data = 12'b111011101110;
20'b00110111010101000111: color_data = 12'b111011101110;
20'b00110111010101001001: color_data = 12'b111011101110;
20'b00110111010101001010: color_data = 12'b111011101110;
20'b00110111010101001011: color_data = 12'b111011101110;
20'b00110111010101001100: color_data = 12'b111011101110;
20'b00110111010101001101: color_data = 12'b111011101110;
20'b00110111010101011111: color_data = 12'b111011101110;
20'b00110111010101100000: color_data = 12'b111011101110;
20'b00110111010101100001: color_data = 12'b111011101110;
20'b00110111010101100010: color_data = 12'b111011101110;
20'b00110111010101100100: color_data = 12'b111111111111;
20'b00110111010101100101: color_data = 12'b111011101110;
20'b00110111010101100110: color_data = 12'b111011101110;
20'b00110111010101100111: color_data = 12'b111011101110;
20'b00110111010101101000: color_data = 12'b111011101110;
20'b00110111010101101111: color_data = 12'b111011101110;
20'b00110111010101110000: color_data = 12'b111011101110;
20'b00110111010101110001: color_data = 12'b111011101110;
20'b00110111010101110010: color_data = 12'b111011101110;
20'b00110111010101110011: color_data = 12'b111111111111;
20'b00110111010101110101: color_data = 12'b111011101110;
20'b00110111010101110110: color_data = 12'b111011101110;
20'b00110111010101110111: color_data = 12'b111011101110;
20'b00110111010101111000: color_data = 12'b111011101110;
20'b00110111010101111001: color_data = 12'b111011101110;
20'b00110111010101111011: color_data = 12'b111011101110;
20'b00110111010101111100: color_data = 12'b111011101110;
20'b00110111010101111101: color_data = 12'b111111111111;
20'b00110111010101111110: color_data = 12'b111011101110;
20'b00110111010110000000: color_data = 12'b111011101110;
20'b00110111010110000001: color_data = 12'b111011101110;
20'b00110111010110000010: color_data = 12'b111011101110;
20'b00110111010110000011: color_data = 12'b111011101110;
20'b00110111010110000100: color_data = 12'b111011101110;
20'b00110111010110000110: color_data = 12'b111011101110;
20'b00110111010110000111: color_data = 12'b111011101110;
20'b00110111010110001000: color_data = 12'b111011101110;
20'b00110111010110001001: color_data = 12'b111011101110;
20'b00110111010110001011: color_data = 12'b111011101110;
20'b00110111010110001100: color_data = 12'b111011101110;
20'b00110111010110001101: color_data = 12'b111011101110;
20'b00110111010110001110: color_data = 12'b111011101110;
20'b00110111010110001111: color_data = 12'b111011101110;
20'b00110111010110010001: color_data = 12'b111011101110;
20'b00110111010110010010: color_data = 12'b111111111111;
20'b00110111010110010011: color_data = 12'b111011101110;
20'b00110111010110010100: color_data = 12'b111011101110;
20'b00110111100011110001: color_data = 12'b111011101110;
20'b00110111100011110010: color_data = 12'b111111111111;
20'b00110111100011110011: color_data = 12'b111011101110;
20'b00110111100011110100: color_data = 12'b111011101110;
20'b00110111100011110101: color_data = 12'b111111111111;
20'b00110111100011110111: color_data = 12'b111011101110;
20'b00110111100011111000: color_data = 12'b111111111111;
20'b00110111100011111001: color_data = 12'b111011101110;
20'b00110111100011111010: color_data = 12'b111111111111;
20'b00110111100011111100: color_data = 12'b111011101110;
20'b00110111100011111101: color_data = 12'b111011101110;
20'b00110111100011111110: color_data = 12'b111011101110;
20'b00110111100011111111: color_data = 12'b111011101110;
20'b00110111100100000001: color_data = 12'b111011101110;
20'b00110111100100000010: color_data = 12'b111111111111;
20'b00110111100100000011: color_data = 12'b111011101110;
20'b00110111100100000100: color_data = 12'b111011101110;
20'b00110111100100000101: color_data = 12'b111111111111;
20'b00110111100100000111: color_data = 12'b111011101110;
20'b00110111100100001000: color_data = 12'b111011101110;
20'b00110111100100001001: color_data = 12'b111111111111;
20'b00110111100100001010: color_data = 12'b111011101110;
20'b00110111100100001011: color_data = 12'b111111111111;
20'b00110111100100010111: color_data = 12'b111011101110;
20'b00110111100100011000: color_data = 12'b111011101110;
20'b00110111100100011001: color_data = 12'b111011101110;
20'b00110111100100011010: color_data = 12'b111011101110;
20'b00110111100100011011: color_data = 12'b111011101110;
20'b00110111100100011101: color_data = 12'b111111111111;
20'b00110111100100011110: color_data = 12'b111011101110;
20'b00110111100100011111: color_data = 12'b111111111111;
20'b00110111100100100000: color_data = 12'b111011101110;
20'b00110111100100100001: color_data = 12'b111111111111;
20'b00110111100100110011: color_data = 12'b111111111111;
20'b00110111100100110100: color_data = 12'b111011101110;
20'b00110111100100110101: color_data = 12'b111111111111;
20'b00110111100100110110: color_data = 12'b111011101110;
20'b00110111100100110111: color_data = 12'b111011101110;
20'b00110111100100111001: color_data = 12'b111011101110;
20'b00110111100100111010: color_data = 12'b111011101110;
20'b00110111100100111011: color_data = 12'b111011101110;
20'b00110111100100111100: color_data = 12'b111011101110;
20'b00110111100101000011: color_data = 12'b111111111111;
20'b00110111100101000100: color_data = 12'b111011101110;
20'b00110111100101000101: color_data = 12'b111111111111;
20'b00110111100101000110: color_data = 12'b111011101110;
20'b00110111100101000111: color_data = 12'b111011101110;
20'b00110111100101001001: color_data = 12'b111011101110;
20'b00110111100101001010: color_data = 12'b111011101110;
20'b00110111100101001011: color_data = 12'b111011101110;
20'b00110111100101001100: color_data = 12'b111011101110;
20'b00110111100101001101: color_data = 12'b111011101110;
20'b00110111100101011111: color_data = 12'b111011101110;
20'b00110111100101100000: color_data = 12'b111111111111;
20'b00110111100101100001: color_data = 12'b111011101110;
20'b00110111100101100010: color_data = 12'b111111111111;
20'b00110111100101100100: color_data = 12'b111011101110;
20'b00110111100101100101: color_data = 12'b111011101110;
20'b00110111100101100110: color_data = 12'b111011101110;
20'b00110111100101100111: color_data = 12'b111011101110;
20'b00110111100101101000: color_data = 12'b111011101110;
20'b00110111100101101111: color_data = 12'b111011101110;
20'b00110111100101110000: color_data = 12'b111011101110;
20'b00110111100101110001: color_data = 12'b111011101110;
20'b00110111100101110010: color_data = 12'b111011101110;
20'b00110111100101110011: color_data = 12'b111011101110;
20'b00110111100101110101: color_data = 12'b111111111111;
20'b00110111100101110110: color_data = 12'b111011101110;
20'b00110111100101110111: color_data = 12'b111111111111;
20'b00110111100101111000: color_data = 12'b111011101110;
20'b00110111100101111001: color_data = 12'b111111111111;
20'b00110111100101111011: color_data = 12'b111011101110;
20'b00110111100101111100: color_data = 12'b111011101110;
20'b00110111100101111101: color_data = 12'b111011101110;
20'b00110111100101111110: color_data = 12'b111011101110;
20'b00110111100110000000: color_data = 12'b111011101110;
20'b00110111100110000001: color_data = 12'b111011101110;
20'b00110111100110000010: color_data = 12'b111011101110;
20'b00110111100110000011: color_data = 12'b111011101110;
20'b00110111100110000100: color_data = 12'b111011101110;
20'b00110111100110000110: color_data = 12'b111111111111;
20'b00110111100110000111: color_data = 12'b111011101110;
20'b00110111100110001000: color_data = 12'b111011101110;
20'b00110111100110001001: color_data = 12'b111111111111;
20'b00110111100110001011: color_data = 12'b111011101110;
20'b00110111100110001100: color_data = 12'b111011101110;
20'b00110111100110001101: color_data = 12'b111011101110;
20'b00110111100110001110: color_data = 12'b111011101110;
20'b00110111100110001111: color_data = 12'b111011101110;
20'b00110111100110010001: color_data = 12'b111011101110;
20'b00110111100110010010: color_data = 12'b111011101110;
20'b00110111100110010011: color_data = 12'b111011101110;
20'b00110111100110010100: color_data = 12'b111011101110;
20'b00110111110011110001: color_data = 12'b111111111111;
20'b00110111110011110010: color_data = 12'b111011101110;
20'b00110111110011110011: color_data = 12'b111011101110;
20'b00110111110011110100: color_data = 12'b111011101110;
20'b00110111110011110101: color_data = 12'b111011101110;
20'b00110111110011110111: color_data = 12'b111011101110;
20'b00110111110011111000: color_data = 12'b111011101110;
20'b00110111110011111001: color_data = 12'b111111111111;
20'b00110111110011111010: color_data = 12'b111011101110;
20'b00110111110011111100: color_data = 12'b111011101110;
20'b00110111110011111101: color_data = 12'b111011101110;
20'b00110111110011111110: color_data = 12'b111011101110;
20'b00110111110011111111: color_data = 12'b111011101110;
20'b00110111110100000001: color_data = 12'b111111111111;
20'b00110111110100000010: color_data = 12'b111011101110;
20'b00110111110100000011: color_data = 12'b111011101110;
20'b00110111110100000100: color_data = 12'b111011101110;
20'b00110111110100000101: color_data = 12'b111011101110;
20'b00110111110100000111: color_data = 12'b111011101110;
20'b00110111110100001000: color_data = 12'b111011101110;
20'b00110111110100001001: color_data = 12'b111011101110;
20'b00110111110100001010: color_data = 12'b111011101110;
20'b00110111110100001011: color_data = 12'b111011101110;
20'b00110111110100010111: color_data = 12'b111011101110;
20'b00110111110100011000: color_data = 12'b111011101110;
20'b00110111110100011001: color_data = 12'b111011101110;
20'b00110111110100011010: color_data = 12'b111011101110;
20'b00110111110100011011: color_data = 12'b111011101110;
20'b00110111110100011101: color_data = 12'b111011101110;
20'b00110111110100011110: color_data = 12'b111111111111;
20'b00110111110100011111: color_data = 12'b111011101110;
20'b00110111110100100000: color_data = 12'b111011101110;
20'b00110111110100100001: color_data = 12'b111011101110;
20'b00110111110100110011: color_data = 12'b111011101110;
20'b00110111110100110100: color_data = 12'b111011101110;
20'b00110111110100110101: color_data = 12'b111011101110;
20'b00110111110100110110: color_data = 12'b111011101110;
20'b00110111110100110111: color_data = 12'b111011101110;
20'b00110111110100111001: color_data = 12'b111111111111;
20'b00110111110100111010: color_data = 12'b111011101110;
20'b00110111110100111011: color_data = 12'b111011101110;
20'b00110111110100111100: color_data = 12'b111011101110;
20'b00110111110101000011: color_data = 12'b111011101110;
20'b00110111110101000100: color_data = 12'b111011101110;
20'b00110111110101000101: color_data = 12'b111011101110;
20'b00110111110101000110: color_data = 12'b111011101110;
20'b00110111110101000111: color_data = 12'b111011101110;
20'b00110111110101001001: color_data = 12'b111011101110;
20'b00110111110101001010: color_data = 12'b111011101110;
20'b00110111110101001011: color_data = 12'b111011101110;
20'b00110111110101001100: color_data = 12'b111011101110;
20'b00110111110101001101: color_data = 12'b111011101110;
20'b00110111110101011111: color_data = 12'b111011101110;
20'b00110111110101100000: color_data = 12'b111011101110;
20'b00110111110101100001: color_data = 12'b111111111111;
20'b00110111110101100010: color_data = 12'b111011101110;
20'b00110111110101100100: color_data = 12'b111011101110;
20'b00110111110101100101: color_data = 12'b111011101110;
20'b00110111110101100110: color_data = 12'b111011101110;
20'b00110111110101100111: color_data = 12'b111011101110;
20'b00110111110101101000: color_data = 12'b111011101110;
20'b00110111110101101111: color_data = 12'b111011101110;
20'b00110111110101110000: color_data = 12'b111011101110;
20'b00110111110101110001: color_data = 12'b111011101110;
20'b00110111110101110010: color_data = 12'b111011101110;
20'b00110111110101110011: color_data = 12'b111011101110;
20'b00110111110101110101: color_data = 12'b111011101110;
20'b00110111110101110110: color_data = 12'b111111111111;
20'b00110111110101110111: color_data = 12'b111011101110;
20'b00110111110101111000: color_data = 12'b111011101110;
20'b00110111110101111001: color_data = 12'b111011101110;
20'b00110111110101111011: color_data = 12'b111011101110;
20'b00110111110101111100: color_data = 12'b111011101110;
20'b00110111110101111101: color_data = 12'b111011101110;
20'b00110111110101111110: color_data = 12'b111011101110;
20'b00110111110110000000: color_data = 12'b111011101110;
20'b00110111110110000001: color_data = 12'b111011101110;
20'b00110111110110000010: color_data = 12'b111011101110;
20'b00110111110110000011: color_data = 12'b111011101110;
20'b00110111110110000100: color_data = 12'b111111111111;
20'b00110111110110000110: color_data = 12'b111011101110;
20'b00110111110110000111: color_data = 12'b111111111111;
20'b00110111110110001000: color_data = 12'b111111111111;
20'b00110111110110001001: color_data = 12'b111011101110;
20'b00110111110110001011: color_data = 12'b111111111111;
20'b00110111110110001100: color_data = 12'b111011101110;
20'b00110111110110001101: color_data = 12'b111011101110;
20'b00110111110110001110: color_data = 12'b111011101110;
20'b00110111110110001111: color_data = 12'b111011101110;
20'b00110111110110010001: color_data = 12'b111111111111;
20'b00110111110110010010: color_data = 12'b111011101110;
20'b00110111110110010011: color_data = 12'b111011101110;
20'b00110111110110010100: color_data = 12'b111011101110;
20'b00111100010011110001: color_data = 12'b000100000001;
20'b00111100010011110010: color_data = 12'b001000000010;
20'b00111100010011110011: color_data = 12'b001000000010;
20'b00111100010011110100: color_data = 12'b001100000010;
20'b00111100010011110101: color_data = 12'b001000000010;
20'b00111100010011110110: color_data = 12'b000100000001;
20'b00111100010011110111: color_data = 12'b000100000001;
20'b00111100010011111000: color_data = 12'b000100000001;
20'b00111100010011111001: color_data = 12'b001000000010;
20'b00111100010011111010: color_data = 12'b000100000001;
20'b00111100010110001010: color_data = 12'b000000000010;
20'b00111100010110001011: color_data = 12'b000000000011;
20'b00111100010110001100: color_data = 12'b000000000010;
20'b00111100010110001101: color_data = 12'b000000000010;
20'b00111100010110001110: color_data = 12'b000000000001;
20'b00111100100011110000: color_data = 12'b001000000010;
20'b00111100100011110001: color_data = 12'b101000111010;
20'b00111100100011110010: color_data = 12'b110000101100;
20'b00111100100011110011: color_data = 12'b110100011101;
20'b00111100100011110100: color_data = 12'b110100011101;
20'b00111100100011110101: color_data = 12'b110100011100;
20'b00111100100011110110: color_data = 12'b010000000100;
20'b00111100100011110111: color_data = 12'b101000111010;
20'b00111100100011111000: color_data = 12'b110000101100;
20'b00111100100011111001: color_data = 12'b110100101100;
20'b00111100100011111010: color_data = 12'b101000111010;
20'b00111100100011111011: color_data = 12'b001000000010;
20'b00111100100011111100: color_data = 12'b000100000000;
20'b00111100100100110010: color_data = 12'b100011111111;
20'b00111100100100110011: color_data = 12'b010111101110;
20'b00111100100100110100: color_data = 12'b011011101111;
20'b00111100100100110101: color_data = 12'b011111101111;
20'b00111100100100110110: color_data = 12'b100011101111;
20'b00111100100100110111: color_data = 12'b000000000001;
20'b00111100100100111000: color_data = 12'b011111101111;
20'b00111100100100111001: color_data = 12'b011011101111;
20'b00111100100100111010: color_data = 12'b010111101111;
20'b00111100100100111011: color_data = 12'b011111101111;
20'b00111100100100111100: color_data = 12'b100111101110;
20'b00111100100110001001: color_data = 12'b000000000010;
20'b00111100100110001010: color_data = 12'b000100101010;
20'b00111100100110001011: color_data = 12'b000000011100;
20'b00111100100110001100: color_data = 12'b000100011101;
20'b00111100100110001101: color_data = 12'b000100011011;
20'b00111100100110001110: color_data = 12'b001000101010;
20'b00111100100110001111: color_data = 12'b000000000011;
20'b00111100100110010000: color_data = 12'b000000000001;
20'b00111100110011101111: color_data = 12'b000100000001;
20'b00111100110011110000: color_data = 12'b001100000011;
20'b00111100110011110001: color_data = 12'b101100101100;
20'b00111100110011110010: color_data = 12'b111000011111;
20'b00111100110011110011: color_data = 12'b111100001111;
20'b00111100110011110100: color_data = 12'b111100001111;
20'b00111100110011110101: color_data = 12'b111100001111;
20'b00111100110011110110: color_data = 12'b010100000101;
20'b00111100110011110111: color_data = 12'b110000101100;
20'b00111100110011111000: color_data = 12'b111100001110;
20'b00111100110011111001: color_data = 12'b111000001110;
20'b00111100110011111010: color_data = 12'b110000101100;
20'b00111100110011111011: color_data = 12'b001100000011;
20'b00111100110011111100: color_data = 12'b000100000001;
20'b00111100110100110010: color_data = 12'b010111101110;
20'b00111100110100110011: color_data = 12'b001111111111;
20'b00111100110100110100: color_data = 12'b001111111111;
20'b00111100110100110101: color_data = 12'b010011101111;
20'b00111100110100110110: color_data = 12'b011011101111;
20'b00111100110100110111: color_data = 12'b000000000001;
20'b00111100110100111000: color_data = 12'b010011101111;
20'b00111100110100111001: color_data = 12'b001111111111;
20'b00111100110100111010: color_data = 12'b001111111111;
20'b00111100110100111011: color_data = 12'b010011101111;
20'b00111100110100111100: color_data = 12'b011111101111;
20'b00111100110100111101: color_data = 12'b000000000001;
20'b00111100110110001001: color_data = 12'b000000000010;
20'b00111100110110001010: color_data = 12'b000000011101;
20'b00111100110110001011: color_data = 12'b000000001111;
20'b00111100110110001100: color_data = 12'b000000001111;
20'b00111100110110001101: color_data = 12'b000000001110;
20'b00111100110110001110: color_data = 12'b001000011011;
20'b00111100110110001111: color_data = 12'b000000000100;
20'b00111100110110010000: color_data = 12'b000000000001;
20'b00111101000011101111: color_data = 12'b000100000001;
20'b00111101000011110000: color_data = 12'b001100000011;
20'b00111101000011110001: color_data = 12'b110000111100;
20'b00111101000011110010: color_data = 12'b110100001110;
20'b00111101000011110011: color_data = 12'b111100001111;
20'b00111101000011110100: color_data = 12'b111100001111;
20'b00111101000011110101: color_data = 12'b111000001110;
20'b00111101000011110110: color_data = 12'b010100000101;
20'b00111101000011110111: color_data = 12'b110000101100;
20'b00111101000011111000: color_data = 12'b111000001110;
20'b00111101000011111001: color_data = 12'b111100011111;
20'b00111101000011111010: color_data = 12'b101100101100;
20'b00111101000011111011: color_data = 12'b001100000011;
20'b00111101000011111100: color_data = 12'b000100000001;
20'b00111101000100100000: color_data = 12'b000000000001;
20'b00111101000100110010: color_data = 12'b010111101110;
20'b00111101000100110011: color_data = 12'b001011111111;
20'b00111101000100110100: color_data = 12'b001011111111;
20'b00111101000100110101: color_data = 12'b001111111111;
20'b00111101000100110110: color_data = 12'b011011101111;
20'b00111101000100110111: color_data = 12'b000000000001;
20'b00111101000100111000: color_data = 12'b010011111111;
20'b00111101000100111001: color_data = 12'b001111101111;
20'b00111101000100111010: color_data = 12'b001111111111;
20'b00111101000100111011: color_data = 12'b010011111111;
20'b00111101000100111100: color_data = 12'b011111111111;
20'b00111101000110001001: color_data = 12'b000000000010;
20'b00111101000110001010: color_data = 12'b000100011101;
20'b00111101000110001011: color_data = 12'b000000001111;
20'b00111101000110001100: color_data = 12'b000000001111;
20'b00111101000110001101: color_data = 12'b000000001110;
20'b00111101000110001110: color_data = 12'b001000101100;
20'b00111101000110001111: color_data = 12'b000000000011;
20'b00111101000110010000: color_data = 12'b000000000001;
20'b00111101010011101111: color_data = 12'b000100000000;
20'b00111101010011110000: color_data = 12'b001100000010;
20'b00111101010011110001: color_data = 12'b101100111011;
20'b00111101010011110010: color_data = 12'b110100011101;
20'b00111101010011110011: color_data = 12'b111000001110;
20'b00111101010011110100: color_data = 12'b111100011111;
20'b00111101010011110101: color_data = 12'b110100011110;
20'b00111101010011110110: color_data = 12'b010100000101;
20'b00111101010011110111: color_data = 12'b101100111011;
20'b00111101010011111000: color_data = 12'b110100011101;
20'b00111101010011111001: color_data = 12'b110100011101;
20'b00111101010011111010: color_data = 12'b101100101011;
20'b00111101010011111011: color_data = 12'b001100000011;
20'b00111101010011111100: color_data = 12'b000100000001;
20'b00111101010100011011: color_data = 12'b000000000001;
20'b00111101010100100000: color_data = 12'b000000000001;
20'b00111101010100100001: color_data = 12'b000000000001;
20'b00111101010100110010: color_data = 12'b011011101110;
20'b00111101010100110011: color_data = 12'b010011111111;
20'b00111101010100110100: color_data = 12'b010011111111;
20'b00111101010100110101: color_data = 12'b010111111111;
20'b00111101010100110110: color_data = 12'b011111101110;
20'b00111101010100110111: color_data = 12'b000000000001;
20'b00111101010100111000: color_data = 12'b010111101111;
20'b00111101010100111001: color_data = 12'b010011101111;
20'b00111101010100111010: color_data = 12'b010011101111;
20'b00111101010100111011: color_data = 12'b010111111111;
20'b00111101010100111100: color_data = 12'b011111101110;
20'b00111101010110001001: color_data = 12'b000000000010;
20'b00111101010110001010: color_data = 12'b000100011011;
20'b00111101010110001011: color_data = 12'b000100001110;
20'b00111101010110001100: color_data = 12'b000000001110;
20'b00111101010110001101: color_data = 12'b000100001101;
20'b00111101010110001110: color_data = 12'b001000101010;
20'b00111101010110001111: color_data = 12'b000000000011;
20'b00111101010110010000: color_data = 12'b000000000001;
20'b00111101010110010001: color_data = 12'b000000000001;
20'b00111101010110010010: color_data = 12'b000000000001;
20'b00111101010110010011: color_data = 12'b000000000001;
20'b00111101100011110000: color_data = 12'b001000000001;
20'b00111101100011110001: color_data = 12'b101001001001;
20'b00111101100011110010: color_data = 12'b101100111011;
20'b00111101100011110011: color_data = 12'b110000101100;
20'b00111101100011110100: color_data = 12'b110000101100;
20'b00111101100011110101: color_data = 12'b110000101100;
20'b00111101100011110110: color_data = 12'b001100000011;
20'b00111101100011110111: color_data = 12'b101001001010;
20'b00111101100011111000: color_data = 12'b101100111011;
20'b00111101100011111001: color_data = 12'b101100111011;
20'b00111101100011111010: color_data = 12'b101001001010;
20'b00111101100011111011: color_data = 12'b001000000010;
20'b00111101100011111100: color_data = 12'b000100000000;
20'b00111101100100010101: color_data = 12'b000000000001;
20'b00111101100100010110: color_data = 12'b000000000001;
20'b00111101100100010111: color_data = 12'b000000000001;
20'b00111101100100011000: color_data = 12'b000000000010;
20'b00111101100100011001: color_data = 12'b000000000010;
20'b00111101100100011010: color_data = 12'b000000000010;
20'b00111101100100011011: color_data = 12'b000000000010;
20'b00111101100100011100: color_data = 12'b000000000001;
20'b00111101100100011101: color_data = 12'b000000000001;
20'b00111101100100011110: color_data = 12'b000000000001;
20'b00111101100100011111: color_data = 12'b000000000010;
20'b00111101100100100000: color_data = 12'b000000000010;
20'b00111101100100100001: color_data = 12'b000000000001;
20'b00111101100100110010: color_data = 12'b000000000001;
20'b00111101100100110011: color_data = 12'b000000000001;
20'b00111101100100110100: color_data = 12'b000000000001;
20'b00111101100100111000: color_data = 12'b000000000001;
20'b00111101100100111001: color_data = 12'b000000000001;
20'b00111101100100111010: color_data = 12'b000000010001;
20'b00111101100101000010: color_data = 12'b000000010000;
20'b00111101100101000011: color_data = 12'b000000010000;
20'b00111101100101000100: color_data = 12'b000000010000;
20'b00111101100101000101: color_data = 12'b000000010000;
20'b00111101100101000110: color_data = 12'b000000010000;
20'b00111101100101000111: color_data = 12'b000000010000;
20'b00111101100101001000: color_data = 12'b000000010000;
20'b00111101100101001001: color_data = 12'b000000010000;
20'b00111101100101001010: color_data = 12'b000000010000;
20'b00111101100101001011: color_data = 12'b000000010000;
20'b00111101100101001100: color_data = 12'b000000010000;
20'b00111101100101001101: color_data = 12'b000000010000;
20'b00111101100101001110: color_data = 12'b000000010000;
20'b00111101100101001111: color_data = 12'b000000010000;
20'b00111101100101010000: color_data = 12'b000000010000;
20'b00111101100101010001: color_data = 12'b000000010000;
20'b00111101100110001001: color_data = 12'b000000000001;
20'b00111101100110001010: color_data = 12'b000000000101;
20'b00111101100110001011: color_data = 12'b000000000110;
20'b00111101100110001100: color_data = 12'b000000000111;
20'b00111101100110001101: color_data = 12'b000000000110;
20'b00111101100110001110: color_data = 12'b000000000100;
20'b00111101100110001111: color_data = 12'b000000000011;
20'b00111101100110010000: color_data = 12'b000000000011;
20'b00111101100110010001: color_data = 12'b000000000011;
20'b00111101100110010010: color_data = 12'b000000000011;
20'b00111101100110010011: color_data = 12'b000000000011;
20'b00111101100110010100: color_data = 12'b000000000001;
20'b00111101110011110000: color_data = 12'b001000000001;
20'b00111101110011110001: color_data = 12'b010000000011;
20'b00111101110011110010: color_data = 12'b010100000100;
20'b00111101110011110011: color_data = 12'b011000000101;
20'b00111101110011110100: color_data = 12'b011000000101;
20'b00111101110011110101: color_data = 12'b010100000101;
20'b00111101110011110110: color_data = 12'b001100000011;
20'b00111101110011110111: color_data = 12'b001000000010;
20'b00111101110011111000: color_data = 12'b001100000010;
20'b00111101110011111001: color_data = 12'b001100000010;
20'b00111101110011111010: color_data = 12'b001000000010;
20'b00111101110011111011: color_data = 12'b000100000001;
20'b00111101110100010110: color_data = 12'b000000000010;
20'b00111101110100010111: color_data = 12'b010110001100;
20'b00111101110100011000: color_data = 12'b001110001100;
20'b00111101110100011001: color_data = 12'b001110001101;
20'b00111101110100011010: color_data = 12'b001110001101;
20'b00111101110100011011: color_data = 12'b010010001101;
20'b00111101110100011100: color_data = 12'b000000000010;
20'b00111101110100011101: color_data = 12'b010110001011;
20'b00111101110100011110: color_data = 12'b010010001100;
20'b00111101110100011111: color_data = 12'b010010001100;
20'b00111101110100100000: color_data = 12'b010110001011;
20'b00111101110100100001: color_data = 12'b000000000001;
20'b00111101110100110010: color_data = 12'b100111101111;
20'b00111101110100110011: color_data = 12'b011111101111;
20'b00111101110100110100: color_data = 12'b011111101111;
20'b00111101110100110101: color_data = 12'b100011101111;
20'b00111101110100110110: color_data = 12'b101011101110;
20'b00111101110100111000: color_data = 12'b100011101110;
20'b00111101110100111001: color_data = 12'b011111101111;
20'b00111101110100111010: color_data = 12'b011111101110;
20'b00111101110100111011: color_data = 12'b100011101110;
20'b00111101110100111100: color_data = 12'b100111101110;
20'b00111101110101000010: color_data = 12'b010111011010;
20'b00111101110101000011: color_data = 12'b010011101001;
20'b00111101110101000100: color_data = 12'b010011101001;
20'b00111101110101000101: color_data = 12'b010111011001;
20'b00111101110101000110: color_data = 12'b011111011010;
20'b00111101110101000111: color_data = 12'b000000010000;
20'b00111101110101001000: color_data = 12'b010011011001;
20'b00111101110101001001: color_data = 12'b010011101001;
20'b00111101110101001010: color_data = 12'b001111101001;
20'b00111101110101001011: color_data = 12'b010111101001;
20'b00111101110101001100: color_data = 12'b011011011001;
20'b00111101110101001101: color_data = 12'b000000010000;
20'b00111101110101001110: color_data = 12'b010111101001;
20'b00111101110101001111: color_data = 12'b010011101001;
20'b00111101110101010000: color_data = 12'b010011101001;
20'b00111101110101010001: color_data = 12'b011011011010;
20'b00111101110110001001: color_data = 12'b000000000001;
20'b00111101110110001010: color_data = 12'b001100101001;
20'b00111101110110001011: color_data = 12'b001000011011;
20'b00111101110110001100: color_data = 12'b000100011100;
20'b00111101110110001101: color_data = 12'b000100011010;
20'b00111101110110001110: color_data = 12'b001000101001;
20'b00111101110110001111: color_data = 12'b000000000100;
20'b00111101110110010000: color_data = 12'b001000101010;
20'b00111101110110010001: color_data = 12'b001000101011;
20'b00111101110110010010: color_data = 12'b001000011011;
20'b00111101110110010011: color_data = 12'b001000101001;
20'b00111101110110010100: color_data = 12'b000000000010;
20'b00111110000011101111: color_data = 12'b000100000000;
20'b00111110000011110000: color_data = 12'b001100000010;
20'b00111110000011110001: color_data = 12'b101100111011;
20'b00111110000011110010: color_data = 12'b110100011101;
20'b00111110000011110011: color_data = 12'b111000001111;
20'b00111110000011110100: color_data = 12'b111000001110;
20'b00111110000011110101: color_data = 12'b110000101100;
20'b00111110000011110110: color_data = 12'b001000000010;
20'b00111110000011111000: color_data = 12'b000100000000;
20'b00111110000011111001: color_data = 12'b000100000001;
20'b00111110000011111010: color_data = 12'b000100000000;
20'b00111110000100010110: color_data = 12'b000000000010;
20'b00111110000100010111: color_data = 12'b010010001101;
20'b00111110000100011000: color_data = 12'b000110001110;
20'b00111110000100011001: color_data = 12'b000010001111;
20'b00111110000100011010: color_data = 12'b000010001111;
20'b00111110000100011011: color_data = 12'b001010001110;
20'b00111110000100011100: color_data = 12'b000000000011;
20'b00111110000100011101: color_data = 12'b010010001100;
20'b00111110000100011110: color_data = 12'b001010001110;
20'b00111110000100011111: color_data = 12'b000110001101;
20'b00111110000100100000: color_data = 12'b010010001100;
20'b00111110000100100001: color_data = 12'b000000000001;
20'b00111110000100110010: color_data = 12'b011011101111;
20'b00111110000100110011: color_data = 12'b010011101111;
20'b00111110000100110100: color_data = 12'b010011101111;
20'b00111110000100110101: color_data = 12'b010111101111;
20'b00111110000100110110: color_data = 12'b100011101111;
20'b00111110000100111000: color_data = 12'b011011101111;
20'b00111110000100111001: color_data = 12'b010111101111;
20'b00111110000100111010: color_data = 12'b010011101111;
20'b00111110000100111011: color_data = 12'b011011101111;
20'b00111110000100111100: color_data = 12'b011111101110;
20'b00111110000101000010: color_data = 12'b010011101001;
20'b00111110000101000011: color_data = 12'b000111111000;
20'b00111110000101000100: color_data = 12'b000111111000;
20'b00111110000101000101: color_data = 12'b001011101001;
20'b00111110000101000110: color_data = 12'b010111101001;
20'b00111110000101000111: color_data = 12'b000000100000;
20'b00111110000101001000: color_data = 12'b001011101000;
20'b00111110000101001001: color_data = 12'b000111111000;
20'b00111110000101001010: color_data = 12'b000111111000;
20'b00111110000101001011: color_data = 12'b001011101001;
20'b00111110000101001100: color_data = 12'b010111101001;
20'b00111110000101001101: color_data = 12'b000000100000;
20'b00111110000101001110: color_data = 12'b001011101000;
20'b00111110000101001111: color_data = 12'b000111111000;
20'b00111110000101010000: color_data = 12'b000111111000;
20'b00111110000101010001: color_data = 12'b010011101001;
20'b00111110000101010010: color_data = 12'b000000010000;
20'b00111110000110001001: color_data = 12'b000000000010;
20'b00111110000110001010: color_data = 12'b000100011011;
20'b00111110000110001011: color_data = 12'b000000001110;
20'b00111110000110001100: color_data = 12'b000000001110;
20'b00111110000110001101: color_data = 12'b000000011101;
20'b00111110000110001110: color_data = 12'b001000101011;
20'b00111110000110001111: color_data = 12'b000000000101;
20'b00111110000110010000: color_data = 12'b000000011100;
20'b00111110000110010001: color_data = 12'b000000001110;
20'b00111110000110010010: color_data = 12'b000000001110;
20'b00111110000110010011: color_data = 12'b000100011011;
20'b00111110000110010100: color_data = 12'b000000000010;
20'b00111110010011101111: color_data = 12'b000100000001;
20'b00111110010011110000: color_data = 12'b001100000011;
20'b00111110010011110001: color_data = 12'b110000101100;
20'b00111110010011110010: color_data = 12'b111000001111;
20'b00111110010011110011: color_data = 12'b111100001111;
20'b00111110010011110100: color_data = 12'b111100001111;
20'b00111110010011110101: color_data = 12'b110100011101;
20'b00111110010011110110: color_data = 12'b001000000010;
20'b00111110010100010110: color_data = 12'b000000000010;
20'b00111110010100010111: color_data = 12'b001110001101;
20'b00111110010100011000: color_data = 12'b000110001111;
20'b00111110010100011001: color_data = 12'b000001111111;
20'b00111110010100011010: color_data = 12'b000001111111;
20'b00111110010100011011: color_data = 12'b000110001110;
20'b00111110010100011100: color_data = 12'b000000000100;
20'b00111110010100011101: color_data = 12'b010010001101;
20'b00111110010100011110: color_data = 12'b000110001111;
20'b00111110010100011111: color_data = 12'b000110001111;
20'b00111110010100100000: color_data = 12'b001110001100;
20'b00111110010100100001: color_data = 12'b000000000001;
20'b00111110010100100010: color_data = 12'b000000000001;
20'b00111110010100110010: color_data = 12'b011011101111;
20'b00111110010100110011: color_data = 12'b001111111111;
20'b00111110010100110100: color_data = 12'b001111101111;
20'b00111110010100110101: color_data = 12'b010011101111;
20'b00111110010100110110: color_data = 12'b011111101111;
20'b00111110010100110111: color_data = 12'b000000000001;
20'b00111110010100111000: color_data = 12'b010011101111;
20'b00111110010100111001: color_data = 12'b001111111111;
20'b00111110010100111010: color_data = 12'b001111111111;
20'b00111110010100111011: color_data = 12'b010011101111;
20'b00111110010100111100: color_data = 12'b011111101111;
20'b00111110010101000010: color_data = 12'b001111111000;
20'b00111110010101000011: color_data = 12'b000011110111;
20'b00111110010101000100: color_data = 12'b000011111000;
20'b00111110010101000101: color_data = 12'b000111111000;
20'b00111110010101000110: color_data = 12'b010011101001;
20'b00111110010101000111: color_data = 12'b000000100000;
20'b00111110010101001000: color_data = 12'b000111111000;
20'b00111110010101001001: color_data = 12'b000011111000;
20'b00111110010101001010: color_data = 12'b000011111000;
20'b00111110010101001011: color_data = 12'b000111111000;
20'b00111110010101001100: color_data = 12'b010011101000;
20'b00111110010101001101: color_data = 12'b000000110000;
20'b00111110010101001110: color_data = 12'b000111111000;
20'b00111110010101001111: color_data = 12'b000011110111;
20'b00111110010101010000: color_data = 12'b000011111000;
20'b00111110010101010001: color_data = 12'b001011111001;
20'b00111110010101010010: color_data = 12'b000000010000;
20'b00111110010110001001: color_data = 12'b000000000011;
20'b00111110010110001010: color_data = 12'b000100011101;
20'b00111110010110001011: color_data = 12'b000000001111;
20'b00111110010110001100: color_data = 12'b000000001111;
20'b00111110010110001101: color_data = 12'b000000011110;
20'b00111110010110001110: color_data = 12'b000100011011;
20'b00111110010110001111: color_data = 12'b000000000110;
20'b00111110010110010000: color_data = 12'b000000001110;
20'b00111110010110010001: color_data = 12'b000000001111;
20'b00111110010110010010: color_data = 12'b000000001111;
20'b00111110010110010011: color_data = 12'b000100011101;
20'b00111110010110010100: color_data = 12'b000000000010;
20'b00111110100011101111: color_data = 12'b000100000001;
20'b00111110100011110000: color_data = 12'b001100000011;
20'b00111110100011110001: color_data = 12'b110000101100;
20'b00111110100011110010: color_data = 12'b111000001110;
20'b00111110100011110011: color_data = 12'b111100001111;
20'b00111110100011110100: color_data = 12'b111100001111;
20'b00111110100011110101: color_data = 12'b110100011101;
20'b00111110100011110110: color_data = 12'b001000000010;
20'b00111110100100010110: color_data = 12'b000000000010;
20'b00111110100100010111: color_data = 12'b010010001101;
20'b00111110100100011000: color_data = 12'b000101111110;
20'b00111110100100011001: color_data = 12'b000010001111;
20'b00111110100100011010: color_data = 12'b000010001111;
20'b00111110100100011011: color_data = 12'b000110001110;
20'b00111110100100011100: color_data = 12'b000000000100;
20'b00111110100100011101: color_data = 12'b001110001101;
20'b00111110100100011110: color_data = 12'b000110001111;
20'b00111110100100011111: color_data = 12'b000010001111;
20'b00111110100100100000: color_data = 12'b010010001101;
20'b00111110100100100001: color_data = 12'b000000000001;
20'b00111110100100110010: color_data = 12'b011011111111;
20'b00111110100100110011: color_data = 12'b001111111111;
20'b00111110100100110100: color_data = 12'b001111111111;
20'b00111110100100110101: color_data = 12'b010011111111;
20'b00111110100100110110: color_data = 12'b011011101111;
20'b00111110100100110111: color_data = 12'b000000000001;
20'b00111110100100111000: color_data = 12'b010111111111;
20'b00111110100100111001: color_data = 12'b010011111111;
20'b00111110100100111010: color_data = 12'b001111111111;
20'b00111110100100111011: color_data = 12'b010011101111;
20'b00111110100100111100: color_data = 12'b011111101110;
20'b00111110100100111101: color_data = 12'b000000010000;
20'b00111110100101000001: color_data = 12'b000000010000;
20'b00111110100101000010: color_data = 12'b001111101000;
20'b00111110100101000011: color_data = 12'b000011110111;
20'b00111110100101000100: color_data = 12'b000011110111;
20'b00111110100101000101: color_data = 12'b000111111000;
20'b00111110100101000110: color_data = 12'b010011101001;
20'b00111110100101000111: color_data = 12'b000000100000;
20'b00111110100101001000: color_data = 12'b000111111000;
20'b00111110100101001001: color_data = 12'b000011110111;
20'b00111110100101001010: color_data = 12'b000011111000;
20'b00111110100101001011: color_data = 12'b000111111000;
20'b00111110100101001100: color_data = 12'b010011101001;
20'b00111110100101001101: color_data = 12'b000000100000;
20'b00111110100101001110: color_data = 12'b000111111000;
20'b00111110100101001111: color_data = 12'b000011110111;
20'b00111110100101010000: color_data = 12'b000011111000;
20'b00111110100101010001: color_data = 12'b001111101001;
20'b00111110100101010010: color_data = 12'b000000010000;
20'b00111110100110001001: color_data = 12'b000000000011;
20'b00111110100110001010: color_data = 12'b000100011101;
20'b00111110100110001011: color_data = 12'b000000001111;
20'b00111110100110001100: color_data = 12'b000000001111;
20'b00111110100110001101: color_data = 12'b000000001101;
20'b00111110100110001110: color_data = 12'b001000011011;
20'b00111110100110001111: color_data = 12'b000000000111;
20'b00111110100110010000: color_data = 12'b000000001110;
20'b00111110100110010001: color_data = 12'b000000001111;
20'b00111110100110010010: color_data = 12'b000000001111;
20'b00111110100110010011: color_data = 12'b001000011101;
20'b00111110100110010100: color_data = 12'b000000000011;
20'b00111110110011110000: color_data = 12'b001000000010;
20'b00111110110011110001: color_data = 12'b101100111011;
20'b00111110110011110010: color_data = 12'b110000101101;
20'b00111110110011110011: color_data = 12'b110000011101;
20'b00111110110011110100: color_data = 12'b110100011110;
20'b00111110110011110101: color_data = 12'b101100101100;
20'b00111110110011110110: color_data = 12'b001000000010;
20'b00111110110100010110: color_data = 12'b000000000001;
20'b00111110110100010111: color_data = 12'b010110001100;
20'b00111110110100011000: color_data = 12'b001110001101;
20'b00111110110100011001: color_data = 12'b001001111101;
20'b00111110110100011010: color_data = 12'b001010001101;
20'b00111110110100011011: color_data = 12'b001110001101;
20'b00111110110100011100: color_data = 12'b000000000011;
20'b00111110110100011101: color_data = 12'b010010001101;
20'b00111110110100011110: color_data = 12'b001001111110;
20'b00111110110100011111: color_data = 12'b001010001110;
20'b00111110110100100000: color_data = 12'b010010001100;
20'b00111110110100100001: color_data = 12'b000000000010;
20'b00111110110100110010: color_data = 12'b011111101110;
20'b00111110110100110011: color_data = 12'b011011101111;
20'b00111110110100110100: color_data = 12'b010111101110;
20'b00111110110100110101: color_data = 12'b011011101110;
20'b00111110110100110110: color_data = 12'b100011101111;
20'b00111110110100110111: color_data = 12'b000000000001;
20'b00111110110100111000: color_data = 12'b011011101111;
20'b00111110110100111001: color_data = 12'b011011101111;
20'b00111110110100111010: color_data = 12'b011011101111;
20'b00111110110100111011: color_data = 12'b011111101111;
20'b00111110110100111100: color_data = 12'b100011101110;
20'b00111110110101000001: color_data = 12'b000000010000;
20'b00111110110101000010: color_data = 12'b001111101000;
20'b00111110110101000011: color_data = 12'b000111111000;
20'b00111110110101000100: color_data = 12'b001011111000;
20'b00111110110101000101: color_data = 12'b001111111000;
20'b00111110110101000110: color_data = 12'b010111101001;
20'b00111110110101000111: color_data = 12'b000000100000;
20'b00111110110101001000: color_data = 12'b010011101001;
20'b00111110110101001001: color_data = 12'b001011101000;
20'b00111110110101001010: color_data = 12'b001111101001;
20'b00111110110101001011: color_data = 12'b010011101001;
20'b00111110110101001100: color_data = 12'b011011011010;
20'b00111110110101001101: color_data = 12'b000000100000;
20'b00111110110101001110: color_data = 12'b001111101000;
20'b00111110110101001111: color_data = 12'b001011111001;
20'b00111110110101010000: color_data = 12'b001011101000;
20'b00111110110101010001: color_data = 12'b010011011001;
20'b00111110110110001001: color_data = 12'b000000000010;
20'b00111110110110001010: color_data = 12'b001000101011;
20'b00111110110110001011: color_data = 12'b000100011100;
20'b00111110110110001100: color_data = 12'b000100011101;
20'b00111110110110001101: color_data = 12'b000100011011;
20'b00111110110110001110: color_data = 12'b001100101001;
20'b00111110110110001111: color_data = 12'b000000000101;
20'b00111110110110010000: color_data = 12'b000100011011;
20'b00111110110110010001: color_data = 12'b000100011101;
20'b00111110110110010010: color_data = 12'b000100011101;
20'b00111110110110010011: color_data = 12'b001000011010;
20'b00111110110110010100: color_data = 12'b000000000010;
20'b00111111000011110000: color_data = 12'b000100000001;
20'b00111111000011110001: color_data = 12'b000100000001;
20'b00111111000011110010: color_data = 12'b000100000010;
20'b00111111000011110011: color_data = 12'b001000000010;
20'b00111111000011110100: color_data = 12'b001000000010;
20'b00111111000011110101: color_data = 12'b000100000001;
20'b00111111000100010111: color_data = 12'b000000000001;
20'b00111111000100011000: color_data = 12'b000000000010;
20'b00111111000100011001: color_data = 12'b000000000001;
20'b00111111000100011010: color_data = 12'b000000000001;
20'b00111111000100011011: color_data = 12'b000000000001;
20'b00111111000100011100: color_data = 12'b000000000001;
20'b00111111000100011101: color_data = 12'b000000000010;
20'b00111111000100011110: color_data = 12'b000000000011;
20'b00111111000100011111: color_data = 12'b000000000011;
20'b00111111000100100000: color_data = 12'b000000000011;
20'b00111111000100100001: color_data = 12'b000000000010;
20'b00111111000101000010: color_data = 12'b000000100000;
20'b00111111000101000011: color_data = 12'b000000100000;
20'b00111111000101000100: color_data = 12'b000000100000;
20'b00111111000101000101: color_data = 12'b000000100000;
20'b00111111000101000110: color_data = 12'b000000010000;
20'b00111111000101000111: color_data = 12'b000000010000;
20'b00111111000101001000: color_data = 12'b000000010000;
20'b00111111000101001001: color_data = 12'b000000010000;
20'b00111111000101001011: color_data = 12'b000000010000;
20'b00111111000101001110: color_data = 12'b000000010000;
20'b00111111000101001111: color_data = 12'b000000010000;
20'b00111111000101010000: color_data = 12'b000000010000;
20'b00111111000101010001: color_data = 12'b000000010000;
20'b00111111000110001001: color_data = 12'b000000000001;
20'b00111111000110001010: color_data = 12'b000000000001;
20'b00111111000110001011: color_data = 12'b000000000010;
20'b00111111000110001100: color_data = 12'b000000000010;
20'b00111111000110001101: color_data = 12'b000000000010;
20'b00111111000110001110: color_data = 12'b000000000010;
20'b00111111000110001111: color_data = 12'b000000000001;
20'b00111111000110010000: color_data = 12'b000000000010;
20'b00111111000110010001: color_data = 12'b000000000010;
20'b00111111000110010010: color_data = 12'b000000000011;
20'b00111111000110010011: color_data = 12'b000000000010;
20'b00111111010011111100: color_data = 12'b111011111110;
20'b00111111010011111101: color_data = 12'b111011111110;
20'b00111111010011111110: color_data = 12'b111011111110;
20'b00111111010011111111: color_data = 12'b111111101110;
20'b00111111010100000000: color_data = 12'b111111101110;
20'b00111111010100000010: color_data = 12'b111011101110;
20'b00111111010100000011: color_data = 12'b111011101110;
20'b00111111010100000100: color_data = 12'b111011101110;
20'b00111111010100000101: color_data = 12'b111011101110;
20'b00111111010100000111: color_data = 12'b111011101110;
20'b00111111010100001000: color_data = 12'b111011101110;
20'b00111111010100001001: color_data = 12'b111011101110;
20'b00111111010100001010: color_data = 12'b111011101110;
20'b00111111010100001011: color_data = 12'b111011101110;
20'b00111111010100011100: color_data = 12'b000000000001;
20'b00111111010100011101: color_data = 12'b011010001011;
20'b00111111010100011110: color_data = 12'b010010001100;
20'b00111111010100011111: color_data = 12'b010010001100;
20'b00111111010100100000: color_data = 12'b010010001100;
20'b00111111010100100001: color_data = 12'b000000000010;
20'b00111111010101000010: color_data = 12'b011011011010;
20'b00111111010101000011: color_data = 12'b001111101000;
20'b00111111010101000100: color_data = 12'b001111101001;
20'b00111111010101000101: color_data = 12'b010011101001;
20'b00111111010101000110: color_data = 12'b011111011011;
20'b00111111010101000111: color_data = 12'b000000010000;
20'b00111111010101010011: color_data = 12'b111111101110;
20'b00111111010101010100: color_data = 12'b111111101110;
20'b00111111010101010101: color_data = 12'b111011101110;
20'b00111111010101010110: color_data = 12'b111011101110;
20'b00111111010101011000: color_data = 12'b111011101110;
20'b00111111010101011001: color_data = 12'b111011111110;
20'b00111111010101011010: color_data = 12'b111011111110;
20'b00111111010101011011: color_data = 12'b111011101110;
20'b00111111010101011100: color_data = 12'b111011101110;
20'b00111111010101011110: color_data = 12'b111011101110;
20'b00111111010101011111: color_data = 12'b111111111111;
20'b00111111010101100000: color_data = 12'b111111111111;
20'b00111111010101100001: color_data = 12'b111011101110;
20'b00111111010101100011: color_data = 12'b111011101110;
20'b00111111010101100100: color_data = 12'b111011101110;
20'b00111111010101100101: color_data = 12'b111011101110;
20'b00111111010101100110: color_data = 12'b111011101110;
20'b00111111010101100111: color_data = 12'b111011101110;
20'b00111111010101110100: color_data = 12'b111011101110;
20'b00111111010101110101: color_data = 12'b111011101110;
20'b00111111010101110110: color_data = 12'b111011101110;
20'b00111111010101110111: color_data = 12'b111011101110;
20'b00111111010101111000: color_data = 12'b111011101110;
20'b00111111010101111010: color_data = 12'b111011101110;
20'b00111111010101111011: color_data = 12'b111011101110;
20'b00111111010101111100: color_data = 12'b111011101110;
20'b00111111010101111101: color_data = 12'b111011101110;
20'b00111111010101111111: color_data = 12'b111011101110;
20'b00111111010110000000: color_data = 12'b111111111111;
20'b00111111010110000001: color_data = 12'b111011101110;
20'b00111111010110000010: color_data = 12'b111011101110;
20'b00111111010110000100: color_data = 12'b111011101110;
20'b00111111010110000101: color_data = 12'b111011101110;
20'b00111111010110000110: color_data = 12'b111011101110;
20'b00111111010110000111: color_data = 12'b111011101110;
20'b00111111010110001000: color_data = 12'b111111101110;
20'b00111111100011111100: color_data = 12'b111011101110;
20'b00111111100011111101: color_data = 12'b111011101110;
20'b00111111100011111110: color_data = 12'b111111101110;
20'b00111111100011111111: color_data = 12'b111011101110;
20'b00111111100100000000: color_data = 12'b111011101110;
20'b00111111100100000010: color_data = 12'b111011101110;
20'b00111111100100000011: color_data = 12'b111011101110;
20'b00111111100100000100: color_data = 12'b111011101110;
20'b00111111100100000101: color_data = 12'b111011101110;
20'b00111111100100000111: color_data = 12'b111011101110;
20'b00111111100100001000: color_data = 12'b111011101110;
20'b00111111100100001001: color_data = 12'b111011101110;
20'b00111111100100001010: color_data = 12'b111011101110;
20'b00111111100100001011: color_data = 12'b111011101110;
20'b00111111100100011100: color_data = 12'b000000000010;
20'b00111111100100011101: color_data = 12'b010010011101;
20'b00111111100100011110: color_data = 12'b000110001110;
20'b00111111100100011111: color_data = 12'b001010001110;
20'b00111111100100100000: color_data = 12'b010010011101;
20'b00111111100100100001: color_data = 12'b000000000010;
20'b00111111100101000001: color_data = 12'b000000010000;
20'b00111111100101000010: color_data = 12'b010011101001;
20'b00111111100101000011: color_data = 12'b001011111000;
20'b00111111100101000100: color_data = 12'b000111111000;
20'b00111111100101000101: color_data = 12'b001011111001;
20'b00111111100101000110: color_data = 12'b010011011001;
20'b00111111100101000111: color_data = 12'b000000010000;
20'b00111111100101010011: color_data = 12'b111111111110;
20'b00111111100101010100: color_data = 12'b111111101110;
20'b00111111100101010101: color_data = 12'b111111101110;
20'b00111111100101010110: color_data = 12'b111011101110;
20'b00111111100101011000: color_data = 12'b111111111111;
20'b00111111100101011001: color_data = 12'b111011101110;
20'b00111111100101011010: color_data = 12'b111111101110;
20'b00111111100101011011: color_data = 12'b111011101110;
20'b00111111100101011100: color_data = 12'b111111111110;
20'b00111111100101011110: color_data = 12'b111011101110;
20'b00111111100101011111: color_data = 12'b111011101110;
20'b00111111100101100000: color_data = 12'b111011101110;
20'b00111111100101100001: color_data = 12'b111011101110;
20'b00111111100101100011: color_data = 12'b111111111111;
20'b00111111100101100100: color_data = 12'b111011101110;
20'b00111111100101100101: color_data = 12'b111011101110;
20'b00111111100101100110: color_data = 12'b111011101110;
20'b00111111100101100111: color_data = 12'b111111111111;
20'b00111111100101110100: color_data = 12'b111011101110;
20'b00111111100101110101: color_data = 12'b111011101110;
20'b00111111100101110110: color_data = 12'b111011101110;
20'b00111111100101110111: color_data = 12'b111011101110;
20'b00111111100101111000: color_data = 12'b111011101110;
20'b00111111100101111010: color_data = 12'b111011101110;
20'b00111111100101111011: color_data = 12'b111011101110;
20'b00111111100101111100: color_data = 12'b111011101110;
20'b00111111100101111101: color_data = 12'b111011101110;
20'b00111111100101111111: color_data = 12'b111011101110;
20'b00111111100110000000: color_data = 12'b111011101110;
20'b00111111100110000001: color_data = 12'b111111111110;
20'b00111111100110000010: color_data = 12'b111011101110;
20'b00111111100110000100: color_data = 12'b111111101111;
20'b00111111100110000101: color_data = 12'b111111111111;
20'b00111111100110000110: color_data = 12'b111011101110;
20'b00111111100110000111: color_data = 12'b111011101110;
20'b00111111100110001000: color_data = 12'b111011101110;
20'b00111111110011111100: color_data = 12'b111011111110;
20'b00111111110011111101: color_data = 12'b111011101110;
20'b00111111110011111110: color_data = 12'b111011101110;
20'b00111111110011111111: color_data = 12'b111111101111;
20'b00111111110100000000: color_data = 12'b111011101110;
20'b00111111110100000010: color_data = 12'b111011101110;
20'b00111111110100000011: color_data = 12'b111011101110;
20'b00111111110100000100: color_data = 12'b111011101110;
20'b00111111110100000101: color_data = 12'b111011101110;
20'b00111111110100000111: color_data = 12'b111011101110;
20'b00111111110100001000: color_data = 12'b111011101110;
20'b00111111110100001001: color_data = 12'b111011101110;
20'b00111111110100001010: color_data = 12'b111011101110;
20'b00111111110100001011: color_data = 12'b111011101110;
20'b00111111110100011100: color_data = 12'b000000000010;
20'b00111111110100011101: color_data = 12'b001010001101;
20'b00111111110100011110: color_data = 12'b000110001111;
20'b00111111110100011111: color_data = 12'b000110001110;
20'b00111111110100100000: color_data = 12'b010010001100;
20'b00111111110100100001: color_data = 12'b000000000010;
20'b00111111110101000001: color_data = 12'b000000010000;
20'b00111111110101000010: color_data = 12'b001111111001;
20'b00111111110101000011: color_data = 12'b000011111000;
20'b00111111110101000100: color_data = 12'b000011110111;
20'b00111111110101000101: color_data = 12'b000111111000;
20'b00111111110101000110: color_data = 12'b010011101001;
20'b00111111110101000111: color_data = 12'b000000010000;
20'b00111111110101010011: color_data = 12'b111011101110;
20'b00111111110101010100: color_data = 12'b111111101110;
20'b00111111110101010101: color_data = 12'b111011101110;
20'b00111111110101010110: color_data = 12'b111011111111;
20'b00111111110101011000: color_data = 12'b111011101110;
20'b00111111110101011001: color_data = 12'b111111101110;
20'b00111111110101011010: color_data = 12'b111111101110;
20'b00111111110101011011: color_data = 12'b111111111110;
20'b00111111110101011100: color_data = 12'b111011101110;
20'b00111111110101011110: color_data = 12'b111011101111;
20'b00111111110101011111: color_data = 12'b111011101110;
20'b00111111110101100000: color_data = 12'b111011101110;
20'b00111111110101100001: color_data = 12'b111011101110;
20'b00111111110101100011: color_data = 12'b111011101110;
20'b00111111110101100100: color_data = 12'b111111111111;
20'b00111111110101100101: color_data = 12'b111011101110;
20'b00111111110101100110: color_data = 12'b111011101110;
20'b00111111110101100111: color_data = 12'b111011101110;
20'b00111111110101110100: color_data = 12'b111011101110;
20'b00111111110101110101: color_data = 12'b111011101110;
20'b00111111110101110110: color_data = 12'b111011101110;
20'b00111111110101110111: color_data = 12'b111011101110;
20'b00111111110101111000: color_data = 12'b111011101110;
20'b00111111110101111010: color_data = 12'b111011101110;
20'b00111111110101111011: color_data = 12'b111011101110;
20'b00111111110101111100: color_data = 12'b111011101110;
20'b00111111110101111101: color_data = 12'b111011101110;
20'b00111111110101111111: color_data = 12'b111011101110;
20'b00111111110110000000: color_data = 12'b111111111110;
20'b00111111110110000001: color_data = 12'b111011101110;
20'b00111111110110000010: color_data = 12'b111011101110;
20'b00111111110110000100: color_data = 12'b111011101110;
20'b00111111110110000101: color_data = 12'b111011101110;
20'b00111111110110000110: color_data = 12'b111011101110;
20'b00111111110110000111: color_data = 12'b111011111110;
20'b00111111110110001000: color_data = 12'b111011101110;
20'b01000000000011111100: color_data = 12'b111011101110;
20'b01000000000011111101: color_data = 12'b111011101110;
20'b01000000000011111110: color_data = 12'b111011101110;
20'b01000000000011111111: color_data = 12'b111011101110;
20'b01000000000100000000: color_data = 12'b111011101110;
20'b01000000000100000010: color_data = 12'b111111111111;
20'b01000000000100000011: color_data = 12'b111011101110;
20'b01000000000100000100: color_data = 12'b111011101110;
20'b01000000000100000101: color_data = 12'b111011101110;
20'b01000000000100000111: color_data = 12'b111011101110;
20'b01000000000100001000: color_data = 12'b111011101110;
20'b01000000000100001001: color_data = 12'b111111111111;
20'b01000000000100001010: color_data = 12'b111011101110;
20'b01000000000100001011: color_data = 12'b111011101110;
20'b01000000000100011011: color_data = 12'b000000000001;
20'b01000000000100011100: color_data = 12'b000000000010;
20'b01000000000100011101: color_data = 12'b001110001110;
20'b01000000000100011110: color_data = 12'b000101111110;
20'b01000000000100011111: color_data = 12'b001010001110;
20'b01000000000100100000: color_data = 12'b010010001100;
20'b01000000000100100001: color_data = 12'b000000000001;
20'b01000000000100100010: color_data = 12'b000000000001;
20'b01000000000101000001: color_data = 12'b000000010000;
20'b01000000000101000010: color_data = 12'b001111101001;
20'b01000000000101000011: color_data = 12'b000011111000;
20'b01000000000101000100: color_data = 12'b000011110111;
20'b01000000000101000101: color_data = 12'b000111111000;
20'b01000000000101000110: color_data = 12'b010111101001;
20'b01000000000101000111: color_data = 12'b000000010000;
20'b01000000000101010011: color_data = 12'b111011101110;
20'b01000000000101010100: color_data = 12'b111011101110;
20'b01000000000101010101: color_data = 12'b111011101110;
20'b01000000000101010110: color_data = 12'b111011101110;
20'b01000000000101011000: color_data = 12'b111011101110;
20'b01000000000101011001: color_data = 12'b111011101110;
20'b01000000000101011010: color_data = 12'b111111101110;
20'b01000000000101011011: color_data = 12'b111111101110;
20'b01000000000101011100: color_data = 12'b111011101110;
20'b01000000000101011110: color_data = 12'b111011101110;
20'b01000000000101011111: color_data = 12'b111011101110;
20'b01000000000101100000: color_data = 12'b111011101110;
20'b01000000000101100001: color_data = 12'b111011101110;
20'b01000000000101100011: color_data = 12'b111011101110;
20'b01000000000101100100: color_data = 12'b111011101110;
20'b01000000000101100101: color_data = 12'b111011101110;
20'b01000000000101100110: color_data = 12'b111011101110;
20'b01000000000101100111: color_data = 12'b111011101110;
20'b01000000000101110100: color_data = 12'b111011101110;
20'b01000000000101110101: color_data = 12'b111011101110;
20'b01000000000101110110: color_data = 12'b111111111111;
20'b01000000000101110111: color_data = 12'b111011101110;
20'b01000000000101111000: color_data = 12'b111011101110;
20'b01000000000101111010: color_data = 12'b111011101110;
20'b01000000000101111011: color_data = 12'b111011101110;
20'b01000000000101111100: color_data = 12'b111011101110;
20'b01000000000101111101: color_data = 12'b111111111111;
20'b01000000000101111111: color_data = 12'b111011101110;
20'b01000000000110000000: color_data = 12'b111011101110;
20'b01000000000110000001: color_data = 12'b111011111110;
20'b01000000000110000010: color_data = 12'b111011101110;
20'b01000000000110000100: color_data = 12'b111011101110;
20'b01000000000110000101: color_data = 12'b111011101110;
20'b01000000000110000110: color_data = 12'b111011101110;
20'b01000000000110000111: color_data = 12'b111011101110;
20'b01000000000110001000: color_data = 12'b111011101110;
20'b01000000010100011100: color_data = 12'b000000000010;
20'b01000000010100011101: color_data = 12'b010010001100;
20'b01000000010100011110: color_data = 12'b001110001101;
20'b01000000010100011111: color_data = 12'b010010001101;
20'b01000000010100100000: color_data = 12'b011010011100;
20'b01000000010100100001: color_data = 12'b000000000001;
20'b01000000010100100010: color_data = 12'b000000000001;
20'b01000000010100100011: color_data = 12'b000000000001;
20'b01000000010101000001: color_data = 12'b000000010000;
20'b01000000010101000010: color_data = 12'b010111101001;
20'b01000000010101000011: color_data = 12'b001111101000;
20'b01000000010101000100: color_data = 12'b001111111000;
20'b01000000010101000101: color_data = 12'b001111101000;
20'b01000000010101000110: color_data = 12'b011011011010;
20'b01000000010101010011: color_data = 12'b111011101110;
20'b01000000010101010100: color_data = 12'b111111111111;
20'b01000000010101010101: color_data = 12'b111011101110;
20'b01000000010101010110: color_data = 12'b111011101110;
20'b01000000010101011000: color_data = 12'b111011101110;
20'b01000000010101011001: color_data = 12'b111111111111;
20'b01000000010101011010: color_data = 12'b111011101110;
20'b01000000010101011011: color_data = 12'b111011101110;
20'b01000000010101011100: color_data = 12'b111011101110;
20'b01000000010101011110: color_data = 12'b111011101110;
20'b01000000010101011111: color_data = 12'b111011101110;
20'b01000000010101100000: color_data = 12'b111011101110;
20'b01000000010101100001: color_data = 12'b111011101110;
20'b01000000010101100011: color_data = 12'b111011101110;
20'b01000000010101100100: color_data = 12'b111011101110;
20'b01000000010101100101: color_data = 12'b111011101110;
20'b01000000010101100110: color_data = 12'b111111111111;
20'b01000000010101100111: color_data = 12'b111011101110;
20'b01000000100011101011: color_data = 12'b111011101110;
20'b01000000100011101100: color_data = 12'b111011101110;
20'b01000000100011101101: color_data = 12'b111011101110;
20'b01000000100011101110: color_data = 12'b111011101110;
20'b01000000100011101111: color_data = 12'b111011101110;
20'b01000000100100000111: color_data = 12'b111011101110;
20'b01000000100100001000: color_data = 12'b111011101110;
20'b01000000100100001001: color_data = 12'b111011101110;
20'b01000000100100001010: color_data = 12'b111011101110;
20'b01000000100100001011: color_data = 12'b111011101110;
20'b01000000100100001101: color_data = 12'b111011101110;
20'b01000000100100001110: color_data = 12'b111011101110;
20'b01000000100100001111: color_data = 12'b111111111111;
20'b01000000100100010000: color_data = 12'b111111101110;
20'b01000000100100010111: color_data = 12'b111111101110;
20'b01000000100100011000: color_data = 12'b111111101110;
20'b01000000100100011001: color_data = 12'b111011101110;
20'b01000000100100011010: color_data = 12'b111011101110;
20'b01000000100100011011: color_data = 12'b111011101111;
20'b01000000100100011101: color_data = 12'b000000000001;
20'b01000000100100011110: color_data = 12'b000000000001;
20'b01000000100100011111: color_data = 12'b000000000001;
20'b01000000100100100000: color_data = 12'b000000000001;
20'b01000000100100100001: color_data = 12'b000000000001;
20'b01000000100100100010: color_data = 12'b000000000001;
20'b01000000100101000011: color_data = 12'b000000010000;
20'b01000000100101000100: color_data = 12'b000000010000;
20'b01000000100101000101: color_data = 12'b000000010000;
20'b01000000100101001000: color_data = 12'b111011101110;
20'b01000000100101001001: color_data = 12'b111011111110;
20'b01000000100101001010: color_data = 12'b111011101110;
20'b01000000100101001011: color_data = 12'b111011111110;
20'b01000000100101001100: color_data = 12'b111011101110;
20'b01000000100101101110: color_data = 12'b111011101110;
20'b01000000100101101111: color_data = 12'b111011101110;
20'b01000000100101110000: color_data = 12'b111111111111;
20'b01000000100101110001: color_data = 12'b111011101110;
20'b01000000100101110010: color_data = 12'b111011101110;
20'b01000000100101110100: color_data = 12'b111011101110;
20'b01000000100101110101: color_data = 12'b111011101110;
20'b01000000100101110110: color_data = 12'b111011101110;
20'b01000000100101110111: color_data = 12'b111011101110;
20'b01000000100101111000: color_data = 12'b111011101110;
20'b01000000110011101011: color_data = 12'b111011101110;
20'b01000000110011101100: color_data = 12'b111011101110;
20'b01000000110011101101: color_data = 12'b111011101110;
20'b01000000110011101110: color_data = 12'b111011101110;
20'b01000000110011101111: color_data = 12'b111011101110;
20'b01000000110100000111: color_data = 12'b111111111111;
20'b01000000110100001000: color_data = 12'b111011101110;
20'b01000000110100001001: color_data = 12'b111011101110;
20'b01000000110100001010: color_data = 12'b111011101110;
20'b01000000110100001011: color_data = 12'b111011101110;
20'b01000000110100001101: color_data = 12'b111011101110;
20'b01000000110100001110: color_data = 12'b111011101110;
20'b01000000110100001111: color_data = 12'b111011101110;
20'b01000000110100010000: color_data = 12'b111011101110;
20'b01000000110100010111: color_data = 12'b111011101110;
20'b01000000110100011000: color_data = 12'b111011101110;
20'b01000000110100011001: color_data = 12'b111011101110;
20'b01000000110100011010: color_data = 12'b111011111111;
20'b01000000110100011011: color_data = 12'b111011101110;
20'b01000000110101001000: color_data = 12'b111111101110;
20'b01000000110101001001: color_data = 12'b111011101110;
20'b01000000110101001010: color_data = 12'b111011101110;
20'b01000000110101001011: color_data = 12'b111011101110;
20'b01000000110101001100: color_data = 12'b111111111110;
20'b01000000110101101110: color_data = 12'b111011101110;
20'b01000000110101101111: color_data = 12'b111011101110;
20'b01000000110101110000: color_data = 12'b111011101110;
20'b01000000110101110001: color_data = 12'b111011101110;
20'b01000000110101110010: color_data = 12'b111011101110;
20'b01000000110101110100: color_data = 12'b111011101110;
20'b01000000110101110101: color_data = 12'b111011101110;
20'b01000000110101110110: color_data = 12'b111011101110;
20'b01000000110101110111: color_data = 12'b111011101110;
20'b01000000110101111000: color_data = 12'b111111111111;
20'b01000001000011101011: color_data = 12'b111011101110;
20'b01000001000011101100: color_data = 12'b111111111111;
20'b01000001000011101101: color_data = 12'b111011101110;
20'b01000001000011101110: color_data = 12'b111011101110;
20'b01000001000011101111: color_data = 12'b111011101110;
20'b01000001000100000111: color_data = 12'b111011101110;
20'b01000001000100001000: color_data = 12'b111011101110;
20'b01000001000100001001: color_data = 12'b111011101110;
20'b01000001000100001010: color_data = 12'b111011101110;
20'b01000001000100001011: color_data = 12'b111011101110;
20'b01000001000100001101: color_data = 12'b111011101110;
20'b01000001000100001110: color_data = 12'b111011101110;
20'b01000001000100001111: color_data = 12'b111011101110;
20'b01000001000100010000: color_data = 12'b111011111111;
20'b01000001000100010111: color_data = 12'b111111111110;
20'b01000001000100011000: color_data = 12'b111111111111;
20'b01000001000100011001: color_data = 12'b111011101110;
20'b01000001000100011010: color_data = 12'b111011101110;
20'b01000001000100011011: color_data = 12'b111011111111;
20'b01000001000101001000: color_data = 12'b111111101110;
20'b01000001000101001001: color_data = 12'b111011101110;
20'b01000001000101001010: color_data = 12'b111011101110;
20'b01000001000101001011: color_data = 12'b111011111110;
20'b01000001000101001100: color_data = 12'b111011101110;
20'b01000001000101101110: color_data = 12'b111011101110;
20'b01000001000101101111: color_data = 12'b111011101110;
20'b01000001000101110000: color_data = 12'b111011101110;
20'b01000001000101110001: color_data = 12'b111011101110;
20'b01000001000101110010: color_data = 12'b111011101110;
20'b01000001000101110100: color_data = 12'b111011101110;
20'b01000001000101110101: color_data = 12'b111011101110;
20'b01000001000101110110: color_data = 12'b111011101110;
20'b01000001000101110111: color_data = 12'b111011101110;
20'b01000001000101111000: color_data = 12'b111011101110;
20'b01000001010011101011: color_data = 12'b111011101110;
20'b01000001010011101100: color_data = 12'b111011101110;
20'b01000001010011101101: color_data = 12'b111011101110;
20'b01000001010011101110: color_data = 12'b111011101110;
20'b01000001010011101111: color_data = 12'b111011101110;
20'b01000001010100000111: color_data = 12'b111011101110;
20'b01000001010100001000: color_data = 12'b111111111111;
20'b01000001010100001001: color_data = 12'b111011101110;
20'b01000001010100001010: color_data = 12'b111011101110;
20'b01000001010100001011: color_data = 12'b111111111111;
20'b01000001010100001101: color_data = 12'b111011101110;
20'b01000001010100001110: color_data = 12'b111111111111;
20'b01000001010100001111: color_data = 12'b111011101110;
20'b01000001010100010000: color_data = 12'b111011101110;
20'b01000001010100010111: color_data = 12'b111011101110;
20'b01000001010100011000: color_data = 12'b111011101110;
20'b01000001010100011001: color_data = 12'b111011101110;
20'b01000001010100011010: color_data = 12'b111011101111;
20'b01000001010100011011: color_data = 12'b111011101111;
20'b01000001010101001000: color_data = 12'b111111101110;
20'b01000001010101001001: color_data = 12'b111011101110;
20'b01000001010101001010: color_data = 12'b111011101110;
20'b01000001010101001011: color_data = 12'b111011101110;
20'b01000001010101001100: color_data = 12'b111011101110;
20'b01000001010101101110: color_data = 12'b111011101110;
20'b01000001010101101111: color_data = 12'b111011101110;
20'b01000001010101110000: color_data = 12'b111011101110;
20'b01000001010101110001: color_data = 12'b111111111111;
20'b01000001010101110010: color_data = 12'b111011101110;
20'b01000001010101110100: color_data = 12'b111111111111;
20'b01000001010101110101: color_data = 12'b111011101110;
20'b01000001010101110110: color_data = 12'b111011101110;
20'b01000001010101110111: color_data = 12'b111111111111;
20'b01000001010101111000: color_data = 12'b111011101110;
20'b01000001100011101011: color_data = 12'b111011101110;
20'b01000001100011101100: color_data = 12'b111011101110;
20'b01000001100011101101: color_data = 12'b111111111111;
20'b01000001100011101110: color_data = 12'b111011101110;
20'b01000001100011101111: color_data = 12'b111011101110;
20'b01000001100100000111: color_data = 12'b111011101110;
20'b01000001100100001000: color_data = 12'b111011101110;
20'b01000001100100001001: color_data = 12'b111011101110;
20'b01000001100100001010: color_data = 12'b111011101110;
20'b01000001100100001011: color_data = 12'b111011101110;
20'b01000001100100001101: color_data = 12'b111111111111;
20'b01000001100100001110: color_data = 12'b111011101110;
20'b01000001100100001111: color_data = 12'b111011101110;
20'b01000001100100010000: color_data = 12'b111011101111;
20'b01000001100100010111: color_data = 12'b111011101110;
20'b01000001100100011000: color_data = 12'b111111101110;
20'b01000001100100011001: color_data = 12'b111011101110;
20'b01000001100100011010: color_data = 12'b111011101111;
20'b01000001100100011011: color_data = 12'b111011101110;
20'b01000001100101001000: color_data = 12'b111111101110;
20'b01000001100101001001: color_data = 12'b111111101110;
20'b01000001100101001010: color_data = 12'b111111101111;
20'b01000001100101001011: color_data = 12'b111011101110;
20'b01000001100101001100: color_data = 12'b111011101111;
20'b01000001100101101110: color_data = 12'b111011101110;
20'b01000001100101101111: color_data = 12'b111011101110;
20'b01000001100101110000: color_data = 12'b111011101110;
20'b01000001100101110001: color_data = 12'b111011101110;
20'b01000001100101110010: color_data = 12'b111111111111;
20'b01000001100101110100: color_data = 12'b111011101110;
20'b01000001100101110101: color_data = 12'b111011101110;
20'b01000001100101110110: color_data = 12'b111011101110;
20'b01000001100101110111: color_data = 12'b111011101110;
20'b01000001100101111000: color_data = 12'b111011101110;
20'b01000010000011101011: color_data = 12'b111011101110;
20'b01000010000011101100: color_data = 12'b111011101110;
20'b01000010000011101101: color_data = 12'b111011101110;
20'b01000010000011101110: color_data = 12'b111011101110;
20'b01000010000011101111: color_data = 12'b111011101110;
20'b01000010000011110001: color_data = 12'b111011101110;
20'b01000010000011110010: color_data = 12'b111011101110;
20'b01000010000011110011: color_data = 12'b111011101110;
20'b01000010000011110100: color_data = 12'b111011101110;
20'b01000010000011110101: color_data = 12'b111011101110;
20'b01000010000100000111: color_data = 12'b111011101110;
20'b01000010000100001000: color_data = 12'b111011101110;
20'b01000010000100001001: color_data = 12'b111011101110;
20'b01000010000100001010: color_data = 12'b111011101110;
20'b01000010000100001011: color_data = 12'b111011101110;
20'b01000010000100001101: color_data = 12'b111011101110;
20'b01000010000100001110: color_data = 12'b111111111111;
20'b01000010000100001111: color_data = 12'b111011101110;
20'b01000010000100010000: color_data = 12'b111011101110;
20'b01000010000100010111: color_data = 12'b111011101110;
20'b01000010000100011000: color_data = 12'b111011101110;
20'b01000010000100011001: color_data = 12'b111011101110;
20'b01000010000100011010: color_data = 12'b111111111110;
20'b01000010000100011011: color_data = 12'b111111101110;
20'b01000010000100011101: color_data = 12'b111111101110;
20'b01000010000100011110: color_data = 12'b111111111111;
20'b01000010000100011111: color_data = 12'b111111101110;
20'b01000010000100100000: color_data = 12'b111111101110;
20'b01000010000100110010: color_data = 12'b111011101110;
20'b01000010000100110011: color_data = 12'b111011101110;
20'b01000010000100110100: color_data = 12'b111011101110;
20'b01000010000100110101: color_data = 12'b111011101110;
20'b01000010000100110110: color_data = 12'b111011101110;
20'b01000010000100111000: color_data = 12'b111011101110;
20'b01000010000100111001: color_data = 12'b111011101110;
20'b01000010000100111010: color_data = 12'b111011101110;
20'b01000010000100111011: color_data = 12'b111011101110;
20'b01000010000100111100: color_data = 12'b111011101110;
20'b01000010000101000010: color_data = 12'b111111101110;
20'b01000010000101000011: color_data = 12'b111111101110;
20'b01000010000101000100: color_data = 12'b111011101110;
20'b01000010000101000101: color_data = 12'b111011111110;
20'b01000010000101000110: color_data = 12'b111011101111;
20'b01000010000101001000: color_data = 12'b111011101111;
20'b01000010000101001001: color_data = 12'b111011101110;
20'b01000010000101001010: color_data = 12'b111011101110;
20'b01000010000101001011: color_data = 12'b111111101110;
20'b01000010000101001100: color_data = 12'b111111111110;
20'b01000010000101101110: color_data = 12'b111011101110;
20'b01000010000101101111: color_data = 12'b111011101110;
20'b01000010000101110000: color_data = 12'b111011101110;
20'b01000010000101110001: color_data = 12'b111111111111;
20'b01000010000101110010: color_data = 12'b111011101110;
20'b01000010000101110100: color_data = 12'b111011101110;
20'b01000010000101110101: color_data = 12'b111011101110;
20'b01000010000101110110: color_data = 12'b111011101110;
20'b01000010000101110111: color_data = 12'b111011101110;
20'b01000010000101111000: color_data = 12'b111011101110;
20'b01000010000110001010: color_data = 12'b111011101110;
20'b01000010000110001011: color_data = 12'b111011101110;
20'b01000010000110001100: color_data = 12'b111111111111;
20'b01000010000110001101: color_data = 12'b111011101110;
20'b01000010000110001110: color_data = 12'b111011101110;
20'b01000010000110010000: color_data = 12'b111011101110;
20'b01000010000110010001: color_data = 12'b111111111111;
20'b01000010000110010010: color_data = 12'b111011101110;
20'b01000010000110010011: color_data = 12'b111011101110;
20'b01000010010011101011: color_data = 12'b111111111111;
20'b01000010010011101100: color_data = 12'b111011101110;
20'b01000010010011101101: color_data = 12'b111111111111;
20'b01000010010011101110: color_data = 12'b111011101110;
20'b01000010010011101111: color_data = 12'b111011101110;
20'b01000010010011110001: color_data = 12'b111011101110;
20'b01000010010011110010: color_data = 12'b111011101110;
20'b01000010010011110011: color_data = 12'b111011101110;
20'b01000010010011110100: color_data = 12'b111011101110;
20'b01000010010011110101: color_data = 12'b111011101110;
20'b01000010010100000111: color_data = 12'b111011101110;
20'b01000010010100001000: color_data = 12'b111011101110;
20'b01000010010100001001: color_data = 12'b111011101110;
20'b01000010010100001010: color_data = 12'b111011101110;
20'b01000010010100001011: color_data = 12'b111011101110;
20'b01000010010100001101: color_data = 12'b111111111111;
20'b01000010010100001110: color_data = 12'b111011101110;
20'b01000010010100001111: color_data = 12'b111111111111;
20'b01000010010100010000: color_data = 12'b111011101110;
20'b01000010010100010111: color_data = 12'b111011101110;
20'b01000010010100011000: color_data = 12'b111011111110;
20'b01000010010100011001: color_data = 12'b111011101110;
20'b01000010010100011010: color_data = 12'b111011101110;
20'b01000010010100011011: color_data = 12'b111011101110;
20'b01000010010100011101: color_data = 12'b111111111110;
20'b01000010010100011110: color_data = 12'b111011101110;
20'b01000010010100011111: color_data = 12'b111111111111;
20'b01000010010100100000: color_data = 12'b111011101110;
20'b01000010010100110010: color_data = 12'b111011101110;
20'b01000010010100110011: color_data = 12'b111011101110;
20'b01000010010100110100: color_data = 12'b111011101110;
20'b01000010010100110101: color_data = 12'b111011101110;
20'b01000010010100110110: color_data = 12'b111011101110;
20'b01000010010100111000: color_data = 12'b111011101110;
20'b01000010010100111001: color_data = 12'b111011101110;
20'b01000010010100111010: color_data = 12'b111111111111;
20'b01000010010100111011: color_data = 12'b111011101110;
20'b01000010010100111100: color_data = 12'b111111111111;
20'b01000010010101000010: color_data = 12'b111111101110;
20'b01000010010101000011: color_data = 12'b111111101110;
20'b01000010010101000100: color_data = 12'b111111101110;
20'b01000010010101000101: color_data = 12'b111011101110;
20'b01000010010101000110: color_data = 12'b111011101111;
20'b01000010010101001000: color_data = 12'b111011101110;
20'b01000010010101001001: color_data = 12'b111011101110;
20'b01000010010101001010: color_data = 12'b111011101110;
20'b01000010010101001011: color_data = 12'b111111111110;
20'b01000010010101001100: color_data = 12'b111011101110;
20'b01000010010101101110: color_data = 12'b111111111111;
20'b01000010010101101111: color_data = 12'b111011101110;
20'b01000010010101110000: color_data = 12'b111111111111;
20'b01000010010101110001: color_data = 12'b111011101110;
20'b01000010010101110010: color_data = 12'b111111111111;
20'b01000010010101110100: color_data = 12'b111011101110;
20'b01000010010101110101: color_data = 12'b111011101110;
20'b01000010010101110110: color_data = 12'b111011101110;
20'b01000010010101110111: color_data = 12'b111011101110;
20'b01000010010101111000: color_data = 12'b111011101110;
20'b01000010010110001010: color_data = 12'b111011101110;
20'b01000010010110001011: color_data = 12'b111111111111;
20'b01000010010110001100: color_data = 12'b111011101110;
20'b01000010010110001101: color_data = 12'b111011101110;
20'b01000010010110001110: color_data = 12'b111111111111;
20'b01000010010110010000: color_data = 12'b111011101110;
20'b01000010010110010001: color_data = 12'b111011101110;
20'b01000010010110010010: color_data = 12'b111011101110;
20'b01000010010110010011: color_data = 12'b111011101110;
20'b01000010100011101011: color_data = 12'b111011101110;
20'b01000010100011101100: color_data = 12'b111111111111;
20'b01000010100011101101: color_data = 12'b111011101110;
20'b01000010100011101110: color_data = 12'b111011101110;
20'b01000010100011101111: color_data = 12'b111011101110;
20'b01000010100011110001: color_data = 12'b111011101110;
20'b01000010100011110010: color_data = 12'b111011101110;
20'b01000010100011110011: color_data = 12'b111011101110;
20'b01000010100011110100: color_data = 12'b111011101110;
20'b01000010100011110101: color_data = 12'b111011101110;
20'b01000010100100000111: color_data = 12'b111011101110;
20'b01000010100100001000: color_data = 12'b111011101110;
20'b01000010100100001001: color_data = 12'b111011101110;
20'b01000010100100001010: color_data = 12'b111011101110;
20'b01000010100100001011: color_data = 12'b111111111111;
20'b01000010100100001101: color_data = 12'b111011101110;
20'b01000010100100001110: color_data = 12'b111011101110;
20'b01000010100100001111: color_data = 12'b111011101110;
20'b01000010100100010000: color_data = 12'b111011101110;
20'b01000010100100010111: color_data = 12'b111011101110;
20'b01000010100100011000: color_data = 12'b111011101110;
20'b01000010100100011001: color_data = 12'b111011101110;
20'b01000010100100011010: color_data = 12'b111011101110;
20'b01000010100100011011: color_data = 12'b111011111111;
20'b01000010100100011101: color_data = 12'b111011101110;
20'b01000010100100011110: color_data = 12'b111011101110;
20'b01000010100100011111: color_data = 12'b111011101110;
20'b01000010100100100000: color_data = 12'b111011101111;
20'b01000010100100110010: color_data = 12'b111011101110;
20'b01000010100100110011: color_data = 12'b111011101110;
20'b01000010100100110100: color_data = 12'b111011101110;
20'b01000010100100110101: color_data = 12'b111011101110;
20'b01000010100100110110: color_data = 12'b111011101110;
20'b01000010100100111000: color_data = 12'b111011101110;
20'b01000010100100111001: color_data = 12'b111011101110;
20'b01000010100100111010: color_data = 12'b111011101110;
20'b01000010100100111011: color_data = 12'b111111111111;
20'b01000010100100111100: color_data = 12'b111011101110;
20'b01000010100101000010: color_data = 12'b111111101111;
20'b01000010100101000011: color_data = 12'b111011101110;
20'b01000010100101000100: color_data = 12'b111011101110;
20'b01000010100101000101: color_data = 12'b111011101111;
20'b01000010100101000110: color_data = 12'b111011101110;
20'b01000010100101001000: color_data = 12'b111011101111;
20'b01000010100101001001: color_data = 12'b111011101110;
20'b01000010100101001010: color_data = 12'b111111101110;
20'b01000010100101001011: color_data = 12'b111111101110;
20'b01000010100101001100: color_data = 12'b111111101110;
20'b01000010100101101110: color_data = 12'b111011101110;
20'b01000010100101101111: color_data = 12'b111011101110;
20'b01000010100101110000: color_data = 12'b111011101110;
20'b01000010100101110001: color_data = 12'b111011101110;
20'b01000010100101110010: color_data = 12'b111011101110;
20'b01000010100101110100: color_data = 12'b111111111111;
20'b01000010100101110101: color_data = 12'b111011101110;
20'b01000010100101110110: color_data = 12'b111011101110;
20'b01000010100101110111: color_data = 12'b111011101110;
20'b01000010100101111000: color_data = 12'b111011101110;
20'b01000010100110001010: color_data = 12'b111111111111;
20'b01000010100110001011: color_data = 12'b111011101110;
20'b01000010100110001100: color_data = 12'b111011101110;
20'b01000010100110001101: color_data = 12'b111011101110;
20'b01000010100110001110: color_data = 12'b111011101110;
20'b01000010100110010000: color_data = 12'b111011101110;
20'b01000010100110010001: color_data = 12'b111011101110;
20'b01000010100110010010: color_data = 12'b111111111111;
20'b01000010100110010011: color_data = 12'b111011101110;
20'b01000010110011101011: color_data = 12'b111011101110;
20'b01000010110011101100: color_data = 12'b111011101110;
20'b01000010110011101101: color_data = 12'b111011101110;
20'b01000010110011101110: color_data = 12'b111011101110;
20'b01000010110011101111: color_data = 12'b111011101110;
20'b01000010110011110001: color_data = 12'b111011101110;
20'b01000010110011110010: color_data = 12'b111011101110;
20'b01000010110011110011: color_data = 12'b111011101110;
20'b01000010110011110100: color_data = 12'b111111111111;
20'b01000010110011110101: color_data = 12'b111011101110;
20'b01000010110100000111: color_data = 12'b111011101110;
20'b01000010110100001000: color_data = 12'b111011101110;
20'b01000010110100001001: color_data = 12'b111011101110;
20'b01000010110100001010: color_data = 12'b111011101110;
20'b01000010110100001011: color_data = 12'b111011101110;
20'b01000010110100001101: color_data = 12'b111111111111;
20'b01000010110100001110: color_data = 12'b111011101110;
20'b01000010110100001111: color_data = 12'b111011101110;
20'b01000010110100010000: color_data = 12'b111011101110;
20'b01000010110100010111: color_data = 12'b111011101110;
20'b01000010110100011000: color_data = 12'b111011101110;
20'b01000010110100011001: color_data = 12'b111011101110;
20'b01000010110100011010: color_data = 12'b111011101110;
20'b01000010110100011011: color_data = 12'b111011101111;
20'b01000010110100011101: color_data = 12'b111011111111;
20'b01000010110100011110: color_data = 12'b111011101110;
20'b01000010110100011111: color_data = 12'b111011101110;
20'b01000010110100100000: color_data = 12'b111011101110;
20'b01000010110100110010: color_data = 12'b111011101110;
20'b01000010110100110011: color_data = 12'b111111111111;
20'b01000010110100110100: color_data = 12'b111011101110;
20'b01000010110100110101: color_data = 12'b111011101110;
20'b01000010110100110110: color_data = 12'b111011101110;
20'b01000010110100111000: color_data = 12'b111011101110;
20'b01000010110100111001: color_data = 12'b111011101110;
20'b01000010110100111010: color_data = 12'b111011101110;
20'b01000010110100111011: color_data = 12'b111011101110;
20'b01000010110100111100: color_data = 12'b111011101110;
20'b01000010110101000010: color_data = 12'b111011101111;
20'b01000010110101000011: color_data = 12'b111111111111;
20'b01000010110101000100: color_data = 12'b111011101110;
20'b01000010110101000101: color_data = 12'b111111101111;
20'b01000010110101000110: color_data = 12'b111011101110;
20'b01000010110101001000: color_data = 12'b111011101110;
20'b01000010110101001001: color_data = 12'b111111101110;
20'b01000010110101001010: color_data = 12'b111111101110;
20'b01000010110101001011: color_data = 12'b111011101110;
20'b01000010110101001100: color_data = 12'b111111111110;
20'b01000010110101101110: color_data = 12'b111011101110;
20'b01000010110101101111: color_data = 12'b111011101110;
20'b01000010110101110000: color_data = 12'b111011101110;
20'b01000010110101110001: color_data = 12'b111011101110;
20'b01000010110101110010: color_data = 12'b111111111111;
20'b01000010110101110100: color_data = 12'b111011101110;
20'b01000010110101110101: color_data = 12'b111011101110;
20'b01000010110101110110: color_data = 12'b111011101110;
20'b01000010110101110111: color_data = 12'b111011101110;
20'b01000010110101111000: color_data = 12'b111011101110;
20'b01000010110110001010: color_data = 12'b111011101110;
20'b01000010110110001011: color_data = 12'b111011101110;
20'b01000010110110001100: color_data = 12'b111011101110;
20'b01000010110110001101: color_data = 12'b111011101110;
20'b01000010110110001110: color_data = 12'b111011101110;
20'b01000010110110010000: color_data = 12'b111011101110;
20'b01000010110110010001: color_data = 12'b111011101110;
20'b01000010110110010010: color_data = 12'b111011101110;
20'b01000010110110010011: color_data = 12'b111011101110;
20'b01000011000011101011: color_data = 12'b111011101110;
20'b01000011000011101100: color_data = 12'b111011101110;
20'b01000011000011101101: color_data = 12'b111011101110;
20'b01000011000011101110: color_data = 12'b111011101110;
20'b01000011000011101111: color_data = 12'b111011101110;
20'b01000011000011110001: color_data = 12'b111111111111;
20'b01000011000011110010: color_data = 12'b111011101110;
20'b01000011000011110011: color_data = 12'b111111111111;
20'b01000011000011110100: color_data = 12'b111011101110;
20'b01000011000011110101: color_data = 12'b111011101110;
20'b01000011000100000111: color_data = 12'b111011101110;
20'b01000011000100001000: color_data = 12'b111011101110;
20'b01000011000100001001: color_data = 12'b111011101110;
20'b01000011000100001010: color_data = 12'b111011101110;
20'b01000011000100001011: color_data = 12'b111011101110;
20'b01000011000100001101: color_data = 12'b111011101110;
20'b01000011000100001110: color_data = 12'b111011101110;
20'b01000011000100001111: color_data = 12'b111011101110;
20'b01000011000100010000: color_data = 12'b111111101111;
20'b01000011000100010111: color_data = 12'b111011101110;
20'b01000011000100011000: color_data = 12'b111011101110;
20'b01000011000100011001: color_data = 12'b111011101110;
20'b01000011000100011010: color_data = 12'b111111101111;
20'b01000011000100011011: color_data = 12'b111111101111;
20'b01000011000100011101: color_data = 12'b111011101110;
20'b01000011000100011110: color_data = 12'b111011101110;
20'b01000011000100011111: color_data = 12'b111011101110;
20'b01000011000100100000: color_data = 12'b111011101110;
20'b01000011000100110010: color_data = 12'b111011101110;
20'b01000011000100110011: color_data = 12'b111011101110;
20'b01000011000100110100: color_data = 12'b111111111111;
20'b01000011000100110101: color_data = 12'b111011101110;
20'b01000011000100110110: color_data = 12'b111111111111;
20'b01000011000100111000: color_data = 12'b111011101110;
20'b01000011000100111001: color_data = 12'b111011101110;
20'b01000011000100111010: color_data = 12'b111011101110;
20'b01000011000100111011: color_data = 12'b111011101110;
20'b01000011000100111100: color_data = 12'b111011101110;
20'b01000011000101000010: color_data = 12'b111011101110;
20'b01000011000101000011: color_data = 12'b111011101110;
20'b01000011000101000100: color_data = 12'b111111111110;
20'b01000011000101000101: color_data = 12'b111011101110;
20'b01000011000101000110: color_data = 12'b111111111110;
20'b01000011000101001000: color_data = 12'b111011101110;
20'b01000011000101001001: color_data = 12'b111011101110;
20'b01000011000101001010: color_data = 12'b111011101110;
20'b01000011000101001011: color_data = 12'b111011101110;
20'b01000011000101001100: color_data = 12'b111011101110;
20'b01000011000101101110: color_data = 12'b111111111111;
20'b01000011000101101111: color_data = 12'b111011101110;
20'b01000011000101110000: color_data = 12'b111011101110;
20'b01000011000101110001: color_data = 12'b111011101110;
20'b01000011000101110010: color_data = 12'b111011101110;
20'b01000011000101110100: color_data = 12'b111011101110;
20'b01000011000101110101: color_data = 12'b111011101110;
20'b01000011000101110110: color_data = 12'b111011101110;
20'b01000011000101110111: color_data = 12'b111011101110;
20'b01000011000101111000: color_data = 12'b111011101110;
20'b01000011000110001010: color_data = 12'b111011101110;
20'b01000011000110001011: color_data = 12'b111011101110;
20'b01000011000110001100: color_data = 12'b111011101110;
20'b01000011000110001101: color_data = 12'b111011101110;
20'b01000011000110001110: color_data = 12'b111011101110;
20'b01000011000110010000: color_data = 12'b111011101110;
20'b01000011000110010001: color_data = 12'b111111111111;
20'b01000011000110010010: color_data = 12'b111011101110;
20'b01000011000110010011: color_data = 12'b111011101110;
20'b01000011100011101011: color_data = 12'b111011101110;
20'b01000011100011101100: color_data = 12'b111011101110;
20'b01000011100011101101: color_data = 12'b111011101110;
20'b01000011100011101110: color_data = 12'b111011101110;
20'b01000011100011101111: color_data = 12'b111011101110;
20'b01000011100011110001: color_data = 12'b111111111111;
20'b01000011100011110010: color_data = 12'b111011101110;
20'b01000011100011110011: color_data = 12'b111011101110;
20'b01000011100011110100: color_data = 12'b111011101110;
20'b01000011100011110101: color_data = 12'b111011101110;
20'b01000011100100000111: color_data = 12'b111011101110;
20'b01000011100100001000: color_data = 12'b111011101110;
20'b01000011100100001001: color_data = 12'b111011101110;
20'b01000011100100001010: color_data = 12'b111011101110;
20'b01000011100100001011: color_data = 12'b111011101110;
20'b01000011100100001101: color_data = 12'b111011101110;
20'b01000011100100001110: color_data = 12'b111011101110;
20'b01000011100100001111: color_data = 12'b111011101110;
20'b01000011100100010000: color_data = 12'b111011101110;
20'b01000011100100010111: color_data = 12'b111011101110;
20'b01000011100100011000: color_data = 12'b111011101110;
20'b01000011100100011001: color_data = 12'b111011101110;
20'b01000011100100011010: color_data = 12'b111011101110;
20'b01000011100100011011: color_data = 12'b111011101110;
20'b01000011100100011101: color_data = 12'b111011101110;
20'b01000011100100011110: color_data = 12'b111011101110;
20'b01000011100100011111: color_data = 12'b111011101110;
20'b01000011100100100000: color_data = 12'b111011101110;
20'b01000011100100110010: color_data = 12'b111011101110;
20'b01000011100100110011: color_data = 12'b111011101110;
20'b01000011100100110100: color_data = 12'b111011101110;
20'b01000011100100110101: color_data = 12'b111011101110;
20'b01000011100100110110: color_data = 12'b111111111111;
20'b01000011100100111000: color_data = 12'b111011101110;
20'b01000011100100111001: color_data = 12'b111011101110;
20'b01000011100100111010: color_data = 12'b111011101110;
20'b01000011100100111011: color_data = 12'b111011101110;
20'b01000011100100111100: color_data = 12'b111011101110;
20'b01000011100101000010: color_data = 12'b111011101110;
20'b01000011100101000011: color_data = 12'b111111101110;
20'b01000011100101000100: color_data = 12'b111011101110;
20'b01000011100101000101: color_data = 12'b111011101110;
20'b01000011100101000110: color_data = 12'b111011111111;
20'b01000011100101001000: color_data = 12'b111011101110;
20'b01000011100101001001: color_data = 12'b111111101110;
20'b01000011100101001010: color_data = 12'b111011101110;
20'b01000011100101001011: color_data = 12'b111111101110;
20'b01000011100101001100: color_data = 12'b111011101110;
20'b01000011100101001110: color_data = 12'b111011101111;
20'b01000011100101001111: color_data = 12'b111011101110;
20'b01000011100101010000: color_data = 12'b111011101110;
20'b01000011100101010001: color_data = 12'b111011101110;
20'b01000011100101010011: color_data = 12'b111011101110;
20'b01000011100101010100: color_data = 12'b111011101110;
20'b01000011100101010101: color_data = 12'b111011101110;
20'b01000011100101010110: color_data = 12'b111111111111;
20'b01000011100101011000: color_data = 12'b111011101110;
20'b01000011100101011001: color_data = 12'b111011101110;
20'b01000011100101011010: color_data = 12'b111011101110;
20'b01000011100101011011: color_data = 12'b111011101110;
20'b01000011100101011100: color_data = 12'b111011101110;
20'b01000011100101101110: color_data = 12'b111011101110;
20'b01000011100101101111: color_data = 12'b111011101110;
20'b01000011100101110000: color_data = 12'b111011101110;
20'b01000011100101110001: color_data = 12'b111011101110;
20'b01000011100101110010: color_data = 12'b111011101110;
20'b01000011100101110100: color_data = 12'b111011101110;
20'b01000011100101110101: color_data = 12'b111011101110;
20'b01000011100101110110: color_data = 12'b111011101110;
20'b01000011100101110111: color_data = 12'b111011101110;
20'b01000011100101111000: color_data = 12'b111011101110;
20'b01000011100101111111: color_data = 12'b111011101110;
20'b01000011100110000000: color_data = 12'b111011101110;
20'b01000011100110000001: color_data = 12'b111011101110;
20'b01000011100110000010: color_data = 12'b111111111111;
20'b01000011100110000100: color_data = 12'b111011101110;
20'b01000011100110000101: color_data = 12'b111011101110;
20'b01000011100110000110: color_data = 12'b111011101110;
20'b01000011100110000111: color_data = 12'b111011101110;
20'b01000011100110001000: color_data = 12'b111111111111;
20'b01000011100110001010: color_data = 12'b111011101110;
20'b01000011100110001011: color_data = 12'b111011101110;
20'b01000011100110001100: color_data = 12'b111011101110;
20'b01000011100110001101: color_data = 12'b111011101110;
20'b01000011100110001110: color_data = 12'b111011101110;
20'b01000011110011101011: color_data = 12'b111011101110;
20'b01000011110011101100: color_data = 12'b111011101110;
20'b01000011110011101101: color_data = 12'b111011101110;
20'b01000011110011101110: color_data = 12'b111011101110;
20'b01000011110011101111: color_data = 12'b111011101110;
20'b01000011110011110001: color_data = 12'b111011101110;
20'b01000011110011110010: color_data = 12'b111011101110;
20'b01000011110011110011: color_data = 12'b111011101110;
20'b01000011110011110100: color_data = 12'b111011101110;
20'b01000011110011110101: color_data = 12'b111011101110;
20'b01000011110100000111: color_data = 12'b111011101110;
20'b01000011110100001000: color_data = 12'b111011101110;
20'b01000011110100001001: color_data = 12'b111011101110;
20'b01000011110100001010: color_data = 12'b111111111111;
20'b01000011110100001011: color_data = 12'b111011101110;
20'b01000011110100001101: color_data = 12'b111011101110;
20'b01000011110100001110: color_data = 12'b111011101110;
20'b01000011110100001111: color_data = 12'b111011101110;
20'b01000011110100010000: color_data = 12'b111011101110;
20'b01000011110100010111: color_data = 12'b111011101110;
20'b01000011110100011000: color_data = 12'b111011101110;
20'b01000011110100011001: color_data = 12'b111011101110;
20'b01000011110100011010: color_data = 12'b111011111110;
20'b01000011110100011011: color_data = 12'b111011101110;
20'b01000011110100011101: color_data = 12'b111011101110;
20'b01000011110100011110: color_data = 12'b111011101110;
20'b01000011110100011111: color_data = 12'b111011101110;
20'b01000011110100100000: color_data = 12'b111011101110;
20'b01000011110100110010: color_data = 12'b111011101110;
20'b01000011110100110011: color_data = 12'b111011101110;
20'b01000011110100110100: color_data = 12'b111011101110;
20'b01000011110100110101: color_data = 12'b111011101110;
20'b01000011110100110110: color_data = 12'b111011101110;
20'b01000011110100111000: color_data = 12'b111011101110;
20'b01000011110100111001: color_data = 12'b111011101110;
20'b01000011110100111010: color_data = 12'b111011101110;
20'b01000011110100111011: color_data = 12'b111011101110;
20'b01000011110100111100: color_data = 12'b111011101110;
20'b01000011110101000010: color_data = 12'b111011101110;
20'b01000011110101000011: color_data = 12'b111011101110;
20'b01000011110101000100: color_data = 12'b111011101110;
20'b01000011110101000101: color_data = 12'b111011101110;
20'b01000011110101000110: color_data = 12'b111011101110;
20'b01000011110101001000: color_data = 12'b111111101110;
20'b01000011110101001001: color_data = 12'b111111101110;
20'b01000011110101001010: color_data = 12'b111011101110;
20'b01000011110101001011: color_data = 12'b111011101110;
20'b01000011110101001100: color_data = 12'b111011101110;
20'b01000011110101001110: color_data = 12'b111111101111;
20'b01000011110101001111: color_data = 12'b111111101111;
20'b01000011110101010000: color_data = 12'b111011101110;
20'b01000011110101010001: color_data = 12'b111011101110;
20'b01000011110101010011: color_data = 12'b111011101110;
20'b01000011110101010100: color_data = 12'b111011101110;
20'b01000011110101010101: color_data = 12'b111011101110;
20'b01000011110101010110: color_data = 12'b111011101110;
20'b01000011110101011000: color_data = 12'b111011101110;
20'b01000011110101011001: color_data = 12'b111011101110;
20'b01000011110101011010: color_data = 12'b111011101110;
20'b01000011110101011011: color_data = 12'b111011101110;
20'b01000011110101011100: color_data = 12'b111011101110;
20'b01000011110101101110: color_data = 12'b111011101110;
20'b01000011110101101111: color_data = 12'b111011101110;
20'b01000011110101110000: color_data = 12'b111011101110;
20'b01000011110101110001: color_data = 12'b111011101110;
20'b01000011110101110010: color_data = 12'b111011101110;
20'b01000011110101110100: color_data = 12'b111011101110;
20'b01000011110101110101: color_data = 12'b111111111111;
20'b01000011110101110110: color_data = 12'b111011101110;
20'b01000011110101110111: color_data = 12'b111011101110;
20'b01000011110101111000: color_data = 12'b111011101110;
20'b01000011110101111111: color_data = 12'b111011101110;
20'b01000011110110000000: color_data = 12'b111011101110;
20'b01000011110110000001: color_data = 12'b111111111111;
20'b01000011110110000010: color_data = 12'b111011101110;
20'b01000011110110000100: color_data = 12'b111011101110;
20'b01000011110110000101: color_data = 12'b111011101110;
20'b01000011110110000110: color_data = 12'b111011101110;
20'b01000011110110000111: color_data = 12'b111011101110;
20'b01000011110110001000: color_data = 12'b111011101110;
20'b01000011110110001010: color_data = 12'b111011101110;
20'b01000011110110001011: color_data = 12'b111011101110;
20'b01000011110110001100: color_data = 12'b111011101110;
20'b01000011110110001101: color_data = 12'b111011101110;
20'b01000011110110001110: color_data = 12'b111011101110;
20'b01000100000011101011: color_data = 12'b111011101110;
20'b01000100000011101100: color_data = 12'b111011101110;
20'b01000100000011101101: color_data = 12'b111011101110;
20'b01000100000011101110: color_data = 12'b111011101110;
20'b01000100000011101111: color_data = 12'b111011101110;
20'b01000100000011110001: color_data = 12'b111011101110;
20'b01000100000011110010: color_data = 12'b111011101110;
20'b01000100000011110011: color_data = 12'b111011101110;
20'b01000100000011110100: color_data = 12'b111011101110;
20'b01000100000011110101: color_data = 12'b111011101110;
20'b01000100000100000111: color_data = 12'b111011101110;
20'b01000100000100001000: color_data = 12'b111011101110;
20'b01000100000100001001: color_data = 12'b111011101110;
20'b01000100000100001010: color_data = 12'b111111111111;
20'b01000100000100001011: color_data = 12'b111011101110;
20'b01000100000100001101: color_data = 12'b111011101110;
20'b01000100000100001110: color_data = 12'b111011101110;
20'b01000100000100001111: color_data = 12'b111011101110;
20'b01000100000100010000: color_data = 12'b111011101110;
20'b01000100000100010111: color_data = 12'b111011101110;
20'b01000100000100011000: color_data = 12'b111011101110;
20'b01000100000100011001: color_data = 12'b111011101110;
20'b01000100000100011010: color_data = 12'b111011101110;
20'b01000100000100011011: color_data = 12'b111011101110;
20'b01000100000100011101: color_data = 12'b111011101110;
20'b01000100000100011110: color_data = 12'b111011101110;
20'b01000100000100011111: color_data = 12'b111011101110;
20'b01000100000100100000: color_data = 12'b111011101110;
20'b01000100000100110010: color_data = 12'b111011101110;
20'b01000100000100110011: color_data = 12'b111011101110;
20'b01000100000100110100: color_data = 12'b111011101110;
20'b01000100000100110101: color_data = 12'b111011101110;
20'b01000100000100110110: color_data = 12'b111011101110;
20'b01000100000100111000: color_data = 12'b111011101110;
20'b01000100000100111001: color_data = 12'b111011101110;
20'b01000100000100111010: color_data = 12'b111011101110;
20'b01000100000100111011: color_data = 12'b111011101110;
20'b01000100000100111100: color_data = 12'b111011101110;
20'b01000100000101000010: color_data = 12'b111011101110;
20'b01000100000101000011: color_data = 12'b111011101110;
20'b01000100000101000100: color_data = 12'b111011101110;
20'b01000100000101000101: color_data = 12'b111011101110;
20'b01000100000101000110: color_data = 12'b111011101110;
20'b01000100000101001000: color_data = 12'b111011101110;
20'b01000100000101001001: color_data = 12'b111111111111;
20'b01000100000101001010: color_data = 12'b111011101110;
20'b01000100000101001011: color_data = 12'b111011101110;
20'b01000100000101001100: color_data = 12'b111111111111;
20'b01000100000101001110: color_data = 12'b111011101110;
20'b01000100000101001111: color_data = 12'b111011101110;
20'b01000100000101010000: color_data = 12'b111011101110;
20'b01000100000101010001: color_data = 12'b111011101110;
20'b01000100000101010011: color_data = 12'b111011101110;
20'b01000100000101010100: color_data = 12'b111011101110;
20'b01000100000101010101: color_data = 12'b111011101110;
20'b01000100000101010110: color_data = 12'b111011101110;
20'b01000100000101011000: color_data = 12'b111011101110;
20'b01000100000101011001: color_data = 12'b111011101110;
20'b01000100000101011010: color_data = 12'b111011101110;
20'b01000100000101011011: color_data = 12'b111011101110;
20'b01000100000101011100: color_data = 12'b111011101110;
20'b01000100000101101110: color_data = 12'b111011101110;
20'b01000100000101101111: color_data = 12'b111011101110;
20'b01000100000101110000: color_data = 12'b111011101110;
20'b01000100000101110001: color_data = 12'b111011101110;
20'b01000100000101110010: color_data = 12'b111011101110;
20'b01000100000101110100: color_data = 12'b111011101110;
20'b01000100000101110101: color_data = 12'b111011101110;
20'b01000100000101110110: color_data = 12'b111011101110;
20'b01000100000101110111: color_data = 12'b111011101110;
20'b01000100000101111000: color_data = 12'b111011101110;
20'b01000100000101111111: color_data = 12'b111011101110;
20'b01000100000110000000: color_data = 12'b111011101110;
20'b01000100000110000001: color_data = 12'b111011101110;
20'b01000100000110000010: color_data = 12'b111011101110;
20'b01000100000110000100: color_data = 12'b111011101110;
20'b01000100000110000101: color_data = 12'b111011101110;
20'b01000100000110000110: color_data = 12'b111111111111;
20'b01000100000110000111: color_data = 12'b111011101110;
20'b01000100000110001000: color_data = 12'b111011101110;
20'b01000100000110001010: color_data = 12'b111011101110;
20'b01000100000110001011: color_data = 12'b111011101110;
20'b01000100000110001100: color_data = 12'b111011101110;
20'b01000100000110001101: color_data = 12'b111111111111;
20'b01000100000110001110: color_data = 12'b111011101110;
20'b01000100010011101011: color_data = 12'b111011101110;
20'b01000100010011101100: color_data = 12'b111011101110;
20'b01000100010011101101: color_data = 12'b111011101110;
20'b01000100010011101110: color_data = 12'b111011101110;
20'b01000100010011101111: color_data = 12'b111011101110;
20'b01000100010011110001: color_data = 12'b111111111111;
20'b01000100010011110010: color_data = 12'b111011101110;
20'b01000100010011110011: color_data = 12'b111011101110;
20'b01000100010011110100: color_data = 12'b111011101110;
20'b01000100010011110101: color_data = 12'b111011101110;
20'b01000100010100000111: color_data = 12'b111011101110;
20'b01000100010100001000: color_data = 12'b111011101110;
20'b01000100010100001001: color_data = 12'b111011101110;
20'b01000100010100001010: color_data = 12'b111011101110;
20'b01000100010100001011: color_data = 12'b111011101110;
20'b01000100010100001101: color_data = 12'b111011101110;
20'b01000100010100001110: color_data = 12'b111011101110;
20'b01000100010100001111: color_data = 12'b111011101110;
20'b01000100010100010000: color_data = 12'b111011101110;
20'b01000100010100010111: color_data = 12'b111011101110;
20'b01000100010100011000: color_data = 12'b111011101110;
20'b01000100010100011001: color_data = 12'b111011101110;
20'b01000100010100011010: color_data = 12'b111011101110;
20'b01000100010100011011: color_data = 12'b111011101110;
20'b01000100010100011101: color_data = 12'b111111111111;
20'b01000100010100011110: color_data = 12'b111011101110;
20'b01000100010100011111: color_data = 12'b111111111111;
20'b01000100010100100000: color_data = 12'b111011101110;
20'b01000100010100110010: color_data = 12'b111011101110;
20'b01000100010100110011: color_data = 12'b111011101110;
20'b01000100010100110100: color_data = 12'b111011101110;
20'b01000100010100110101: color_data = 12'b111011101110;
20'b01000100010100110110: color_data = 12'b111011101110;
20'b01000100010100111000: color_data = 12'b111011101110;
20'b01000100010100111001: color_data = 12'b111111111111;
20'b01000100010100111010: color_data = 12'b111011101110;
20'b01000100010100111011: color_data = 12'b111011101110;
20'b01000100010100111100: color_data = 12'b111011101110;
20'b01000100010101000010: color_data = 12'b111011101110;
20'b01000100010101000011: color_data = 12'b111011101110;
20'b01000100010101000100: color_data = 12'b111011101110;
20'b01000100010101000101: color_data = 12'b111011101110;
20'b01000100010101000110: color_data = 12'b111011101110;
20'b01000100010101001000: color_data = 12'b111011101110;
20'b01000100010101001001: color_data = 12'b111011101110;
20'b01000100010101001010: color_data = 12'b111111111111;
20'b01000100010101001011: color_data = 12'b111011101110;
20'b01000100010101001100: color_data = 12'b111011101110;
20'b01000100010101001110: color_data = 12'b111111111111;
20'b01000100010101001111: color_data = 12'b111011101110;
20'b01000100010101010000: color_data = 12'b111011101110;
20'b01000100010101010001: color_data = 12'b111011101110;
20'b01000100010101010011: color_data = 12'b111011101110;
20'b01000100010101010100: color_data = 12'b111011101110;
20'b01000100010101010101: color_data = 12'b111011101110;
20'b01000100010101010110: color_data = 12'b111111111111;
20'b01000100010101011000: color_data = 12'b111011101110;
20'b01000100010101011001: color_data = 12'b111011101110;
20'b01000100010101011010: color_data = 12'b111011101110;
20'b01000100010101011011: color_data = 12'b111011101110;
20'b01000100010101011100: color_data = 12'b111011101110;
20'b01000100010101101110: color_data = 12'b111011101110;
20'b01000100010101101111: color_data = 12'b111011101110;
20'b01000100010101110000: color_data = 12'b111111111111;
20'b01000100010101110001: color_data = 12'b111011101110;
20'b01000100010101110010: color_data = 12'b111111111111;
20'b01000100010101110100: color_data = 12'b111011101110;
20'b01000100010101110101: color_data = 12'b111011101110;
20'b01000100010101110110: color_data = 12'b111011101110;
20'b01000100010101110111: color_data = 12'b111011101110;
20'b01000100010101111000: color_data = 12'b111011101110;
20'b01000100010101111111: color_data = 12'b111011101110;
20'b01000100010110000000: color_data = 12'b111011101110;
20'b01000100010110000001: color_data = 12'b111011101110;
20'b01000100010110000010: color_data = 12'b111011101110;
20'b01000100010110000100: color_data = 12'b111011101110;
20'b01000100010110000101: color_data = 12'b111011101110;
20'b01000100010110000110: color_data = 12'b111011101110;
20'b01000100010110000111: color_data = 12'b111111111111;
20'b01000100010110001000: color_data = 12'b111011101110;
20'b01000100010110001010: color_data = 12'b111111111111;
20'b01000100010110001011: color_data = 12'b111011101110;
20'b01000100010110001100: color_data = 12'b111011101110;
20'b01000100010110001101: color_data = 12'b111111111111;
20'b01000100010110001110: color_data = 12'b111011101110;
20'b01000100110011101011: color_data = 12'b111011101110;
20'b01000100110011101100: color_data = 12'b111011101110;
20'b01000100110011101101: color_data = 12'b111011101110;
20'b01000100110011101110: color_data = 12'b111011101110;
20'b01000100110011101111: color_data = 12'b111011101110;
20'b01000100110011110001: color_data = 12'b111111111111;
20'b01000100110011110010: color_data = 12'b111011101110;
20'b01000100110011110011: color_data = 12'b111111111111;
20'b01000100110011110100: color_data = 12'b111011101110;
20'b01000100110011110101: color_data = 12'b111011101110;
20'b01000100110100000111: color_data = 12'b111011101110;
20'b01000100110100001000: color_data = 12'b111011101110;
20'b01000100110100001001: color_data = 12'b111011101110;
20'b01000100110100001010: color_data = 12'b111011101110;
20'b01000100110100001011: color_data = 12'b111011101110;
20'b01000100110100001101: color_data = 12'b111011101110;
20'b01000100110100001110: color_data = 12'b111011101110;
20'b01000100110100001111: color_data = 12'b111011101110;
20'b01000100110100010000: color_data = 12'b111011101110;
20'b01000100110100010111: color_data = 12'b111011101110;
20'b01000100110100011000: color_data = 12'b111011101110;
20'b01000100110100011001: color_data = 12'b111011101110;
20'b01000100110100011010: color_data = 12'b111011101110;
20'b01000100110100011011: color_data = 12'b111011101110;
20'b01000100110100011101: color_data = 12'b111011101110;
20'b01000100110100011110: color_data = 12'b111011101110;
20'b01000100110100011111: color_data = 12'b111011101110;
20'b01000100110100100000: color_data = 12'b111011101110;
20'b01000100110100110010: color_data = 12'b111011101110;
20'b01000100110100110011: color_data = 12'b111011101110;
20'b01000100110100110100: color_data = 12'b111011101110;
20'b01000100110100110101: color_data = 12'b111011101110;
20'b01000100110100110110: color_data = 12'b111011101110;
20'b01000100110100111000: color_data = 12'b111011101110;
20'b01000100110100111001: color_data = 12'b111011101110;
20'b01000100110100111010: color_data = 12'b111111111111;
20'b01000100110100111011: color_data = 12'b111011101110;
20'b01000100110100111100: color_data = 12'b111011101110;
20'b01000100110101000010: color_data = 12'b111011101110;
20'b01000100110101000011: color_data = 12'b111011101110;
20'b01000100110101000100: color_data = 12'b111011101110;
20'b01000100110101000101: color_data = 12'b111011101110;
20'b01000100110101000110: color_data = 12'b111011101110;
20'b01000100110101001000: color_data = 12'b111011101110;
20'b01000100110101001001: color_data = 12'b111011101110;
20'b01000100110101001010: color_data = 12'b111011101110;
20'b01000100110101001011: color_data = 12'b111011101110;
20'b01000100110101001100: color_data = 12'b111011101110;
20'b01000100110101101110: color_data = 12'b111111111111;
20'b01000100110101101111: color_data = 12'b111011101110;
20'b01000100110101110000: color_data = 12'b111011101110;
20'b01000100110101110001: color_data = 12'b111011101110;
20'b01000100110101110010: color_data = 12'b111011101110;
20'b01000100110101110100: color_data = 12'b111011101110;
20'b01000100110101110101: color_data = 12'b111011101110;
20'b01000100110101110110: color_data = 12'b111011101110;
20'b01000100110101110111: color_data = 12'b111011101110;
20'b01000100110101111000: color_data = 12'b111011101110;
20'b01000100110101111010: color_data = 12'b111011101110;
20'b01000100110101111011: color_data = 12'b111011101110;
20'b01000100110101111100: color_data = 12'b111011101110;
20'b01000100110101111101: color_data = 12'b111011101110;
20'b01000100110101111111: color_data = 12'b111011101110;
20'b01000100110110000000: color_data = 12'b111011101110;
20'b01000100110110000001: color_data = 12'b111011101110;
20'b01000100110110000010: color_data = 12'b111011101110;
20'b01000101000011101011: color_data = 12'b111011101110;
20'b01000101000011101100: color_data = 12'b111011101110;
20'b01000101000011101101: color_data = 12'b111011101110;
20'b01000101000011101110: color_data = 12'b111011101110;
20'b01000101000011101111: color_data = 12'b111011101110;
20'b01000101000011110001: color_data = 12'b111011101110;
20'b01000101000011110010: color_data = 12'b111011101110;
20'b01000101000011110011: color_data = 12'b111011101110;
20'b01000101000011110100: color_data = 12'b111111111111;
20'b01000101000011110101: color_data = 12'b111011101110;
20'b01000101000100000111: color_data = 12'b111011101110;
20'b01000101000100001000: color_data = 12'b111011101110;
20'b01000101000100001001: color_data = 12'b111011101110;
20'b01000101000100001010: color_data = 12'b111011101110;
20'b01000101000100001011: color_data = 12'b111011101110;
20'b01000101000100001101: color_data = 12'b111111111111;
20'b01000101000100001110: color_data = 12'b111011101110;
20'b01000101000100001111: color_data = 12'b111011101110;
20'b01000101000100010000: color_data = 12'b111011101110;
20'b01000101000100010111: color_data = 12'b111011101110;
20'b01000101000100011000: color_data = 12'b111011101110;
20'b01000101000100011001: color_data = 12'b111111111111;
20'b01000101000100011010: color_data = 12'b111111111111;
20'b01000101000100011011: color_data = 12'b111011101110;
20'b01000101000100011101: color_data = 12'b111011101110;
20'b01000101000100011110: color_data = 12'b111011101110;
20'b01000101000100011111: color_data = 12'b111011101110;
20'b01000101000100100000: color_data = 12'b111111111111;
20'b01000101000100110010: color_data = 12'b111011101110;
20'b01000101000100110011: color_data = 12'b111011101110;
20'b01000101000100110100: color_data = 12'b111011101110;
20'b01000101000100110101: color_data = 12'b111111111111;
20'b01000101000100110110: color_data = 12'b111011101110;
20'b01000101000100111000: color_data = 12'b111011101110;
20'b01000101000100111001: color_data = 12'b111011101110;
20'b01000101000100111010: color_data = 12'b111011101110;
20'b01000101000100111011: color_data = 12'b111011101110;
20'b01000101000100111100: color_data = 12'b111111111111;
20'b01000101000101000010: color_data = 12'b111011101110;
20'b01000101000101000011: color_data = 12'b111011101110;
20'b01000101000101000100: color_data = 12'b111011101110;
20'b01000101000101000101: color_data = 12'b111111111111;
20'b01000101000101000110: color_data = 12'b111011101110;
20'b01000101000101001000: color_data = 12'b111111111111;
20'b01000101000101001001: color_data = 12'b111011101110;
20'b01000101000101001010: color_data = 12'b111011101110;
20'b01000101000101001011: color_data = 12'b111011101110;
20'b01000101000101001100: color_data = 12'b111011101110;
20'b01000101000101101110: color_data = 12'b111011101110;
20'b01000101000101101111: color_data = 12'b111111111111;
20'b01000101000101110000: color_data = 12'b111011101110;
20'b01000101000101110001: color_data = 12'b111011101110;
20'b01000101000101110010: color_data = 12'b111011101110;
20'b01000101000101110100: color_data = 12'b111011101110;
20'b01000101000101110101: color_data = 12'b111111111111;
20'b01000101000101110110: color_data = 12'b111111111111;
20'b01000101000101110111: color_data = 12'b111011101110;
20'b01000101000101111000: color_data = 12'b111011101110;
20'b01000101000101111010: color_data = 12'b111011101110;
20'b01000101000101111011: color_data = 12'b111011101110;
20'b01000101000101111100: color_data = 12'b111011101110;
20'b01000101000101111101: color_data = 12'b111011101110;
20'b01000101000101111111: color_data = 12'b111011101110;
20'b01000101000110000000: color_data = 12'b111011101110;
20'b01000101000110000001: color_data = 12'b111111111111;
20'b01000101000110000010: color_data = 12'b111011101110;
20'b01000101010011101011: color_data = 12'b111011101110;
20'b01000101010011101100: color_data = 12'b111111111111;
20'b01000101010011101101: color_data = 12'b111011101110;
20'b01000101010011101110: color_data = 12'b111011101110;
20'b01000101010011101111: color_data = 12'b111011101110;
20'b01000101010011110001: color_data = 12'b111011101110;
20'b01000101010011110010: color_data = 12'b111011101110;
20'b01000101010011110011: color_data = 12'b111011101110;
20'b01000101010011110100: color_data = 12'b111011101110;
20'b01000101010011110101: color_data = 12'b111011101110;
20'b01000101010100000111: color_data = 12'b111011101110;
20'b01000101010100001000: color_data = 12'b111011101110;
20'b01000101010100001001: color_data = 12'b111011101110;
20'b01000101010100001010: color_data = 12'b111011101110;
20'b01000101010100001011: color_data = 12'b111111111111;
20'b01000101010100001101: color_data = 12'b111011101110;
20'b01000101010100001110: color_data = 12'b111011101110;
20'b01000101010100001111: color_data = 12'b111011101110;
20'b01000101010100010000: color_data = 12'b111011101110;
20'b01000101010100010111: color_data = 12'b111011101110;
20'b01000101010100011000: color_data = 12'b111011101110;
20'b01000101010100011001: color_data = 12'b111011101110;
20'b01000101010100011010: color_data = 12'b111011101110;
20'b01000101010100011011: color_data = 12'b111011101110;
20'b01000101010100011101: color_data = 12'b111011101110;
20'b01000101010100011110: color_data = 12'b111111111111;
20'b01000101010100011111: color_data = 12'b111011101110;
20'b01000101010100100000: color_data = 12'b111011101110;
20'b01000101010100110010: color_data = 12'b111011101110;
20'b01000101010100110011: color_data = 12'b111111111111;
20'b01000101010100110100: color_data = 12'b111111111111;
20'b01000101010100110101: color_data = 12'b111011101110;
20'b01000101010100110110: color_data = 12'b111011101110;
20'b01000101010100111000: color_data = 12'b111011101110;
20'b01000101010100111001: color_data = 12'b111011101110;
20'b01000101010100111010: color_data = 12'b111011101110;
20'b01000101010100111011: color_data = 12'b111011101110;
20'b01000101010100111100: color_data = 12'b111011101110;
20'b01000101010101000010: color_data = 12'b111011101110;
20'b01000101010101000011: color_data = 12'b111111111111;
20'b01000101010101000100: color_data = 12'b111111111111;
20'b01000101010101000101: color_data = 12'b111011101110;
20'b01000101010101000110: color_data = 12'b111011101110;
20'b01000101010101001000: color_data = 12'b111011101110;
20'b01000101010101001001: color_data = 12'b111111111111;
20'b01000101010101001010: color_data = 12'b111011101110;
20'b01000101010101001011: color_data = 12'b111011101110;
20'b01000101010101001100: color_data = 12'b111011101110;
20'b01000101010101101110: color_data = 12'b111011101110;
20'b01000101010101101111: color_data = 12'b111011101110;
20'b01000101010101110000: color_data = 12'b111011101110;
20'b01000101010101110001: color_data = 12'b111111111111;
20'b01000101010101110010: color_data = 12'b111011101110;
20'b01000101010101110100: color_data = 12'b111011101110;
20'b01000101010101110101: color_data = 12'b111011101110;
20'b01000101010101110110: color_data = 12'b111011101110;
20'b01000101010101110111: color_data = 12'b111011101110;
20'b01000101010101111000: color_data = 12'b111011101110;
20'b01000101010101111010: color_data = 12'b111011101110;
20'b01000101010101111011: color_data = 12'b111011101110;
20'b01000101010101111100: color_data = 12'b111011101110;
20'b01000101010101111101: color_data = 12'b111011101110;
20'b01000101010101111111: color_data = 12'b111011101110;
20'b01000101010110000000: color_data = 12'b111011101110;
20'b01000101010110000001: color_data = 12'b111011101110;
20'b01000101010110000010: color_data = 12'b111011101110;
20'b01000101100011101011: color_data = 12'b111111111111;
20'b01000101100011101100: color_data = 12'b111011101110;
20'b01000101100011101101: color_data = 12'b111111111111;
20'b01000101100011101110: color_data = 12'b111011101110;
20'b01000101100011101111: color_data = 12'b111011101110;
20'b01000101100011110001: color_data = 12'b111011101110;
20'b01000101100011110010: color_data = 12'b111011101110;
20'b01000101100011110011: color_data = 12'b111011101110;
20'b01000101100011110100: color_data = 12'b111011101110;
20'b01000101100011110101: color_data = 12'b111011101110;
20'b01000101100100000111: color_data = 12'b111011101110;
20'b01000101100100001000: color_data = 12'b111011101110;
20'b01000101100100001001: color_data = 12'b111011101110;
20'b01000101100100001010: color_data = 12'b111011101110;
20'b01000101100100001011: color_data = 12'b111011101110;
20'b01000101100100001101: color_data = 12'b111111111111;
20'b01000101100100001110: color_data = 12'b111011101110;
20'b01000101100100001111: color_data = 12'b111111111111;
20'b01000101100100010000: color_data = 12'b111111111111;
20'b01000101100100010111: color_data = 12'b111011101110;
20'b01000101100100011000: color_data = 12'b111111111111;
20'b01000101100100011001: color_data = 12'b111111111111;
20'b01000101100100011010: color_data = 12'b111011101110;
20'b01000101100100011011: color_data = 12'b111011101110;
20'b01000101100100011101: color_data = 12'b111011101110;
20'b01000101100100011110: color_data = 12'b111011101110;
20'b01000101100100011111: color_data = 12'b111011101110;
20'b01000101100100100000: color_data = 12'b111011101110;
20'b01000101100100110010: color_data = 12'b111111111111;
20'b01000101100100110011: color_data = 12'b111011101110;
20'b01000101100100110100: color_data = 12'b111011101110;
20'b01000101100100110101: color_data = 12'b111011101110;
20'b01000101100100110110: color_data = 12'b111011101110;
20'b01000101100100111000: color_data = 12'b111011101110;
20'b01000101100100111001: color_data = 12'b111011101110;
20'b01000101100100111010: color_data = 12'b111011101110;
20'b01000101100100111011: color_data = 12'b111011101110;
20'b01000101100100111100: color_data = 12'b111011101110;
20'b01000101100101000010: color_data = 12'b111111111111;
20'b01000101100101000011: color_data = 12'b111011101110;
20'b01000101100101000100: color_data = 12'b111011101110;
20'b01000101100101000101: color_data = 12'b111011101110;
20'b01000101100101000110: color_data = 12'b111011101110;
20'b01000101100101001000: color_data = 12'b111011101110;
20'b01000101100101001001: color_data = 12'b111011101110;
20'b01000101100101001010: color_data = 12'b111011101110;
20'b01000101100101001011: color_data = 12'b111011101110;
20'b01000101100101001100: color_data = 12'b111011101110;
20'b01000101100101101110: color_data = 12'b111111111111;
20'b01000101100101101111: color_data = 12'b111011101110;
20'b01000101100101110000: color_data = 12'b111011101110;
20'b01000101100101110001: color_data = 12'b111011101110;
20'b01000101100101110010: color_data = 12'b111011101110;
20'b01000101100101110100: color_data = 12'b111011101110;
20'b01000101100101110101: color_data = 12'b111011101110;
20'b01000101100101110110: color_data = 12'b111111111111;
20'b01000101100101110111: color_data = 12'b111111111111;
20'b01000101100101111000: color_data = 12'b111011101110;
20'b01000101100101111010: color_data = 12'b111111111111;
20'b01000101100101111011: color_data = 12'b111011101110;
20'b01000101100101111100: color_data = 12'b111011101110;
20'b01000101100101111101: color_data = 12'b111111111111;
20'b01000101100101111111: color_data = 12'b111011101110;
20'b01000101100110000000: color_data = 12'b111011101110;
20'b01000101100110000001: color_data = 12'b111011101110;
20'b01000101100110000010: color_data = 12'b111011101110;
20'b01000101110011101011: color_data = 12'b111011101110;
20'b01000101110011101100: color_data = 12'b111011101110;
20'b01000101110011101101: color_data = 12'b111011101110;
20'b01000101110011101110: color_data = 12'b111011101110;
20'b01000101110011101111: color_data = 12'b111011101110;
20'b01000101110011110001: color_data = 12'b111011101110;
20'b01000101110011110010: color_data = 12'b111011101110;
20'b01000101110011110011: color_data = 12'b111011101110;
20'b01000101110011110100: color_data = 12'b111011101110;
20'b01000101110011110101: color_data = 12'b111011101110;
20'b01000101110100000111: color_data = 12'b111011101110;
20'b01000101110100001000: color_data = 12'b111011101110;
20'b01000101110100001001: color_data = 12'b111011101110;
20'b01000101110100001010: color_data = 12'b111011101110;
20'b01000101110100001011: color_data = 12'b111011101110;
20'b01000101110100001101: color_data = 12'b111011101110;
20'b01000101110100001110: color_data = 12'b111111111111;
20'b01000101110100001111: color_data = 12'b111011101110;
20'b01000101110100010000: color_data = 12'b111011101110;
20'b01000110000100010111: color_data = 12'b111011101110;
20'b01000110000100011000: color_data = 12'b111011101110;
20'b01000110000100011001: color_data = 12'b111011101110;
20'b01000110000100011010: color_data = 12'b111011101110;
20'b01000110000100011011: color_data = 12'b111011101110;
20'b01000110000100011101: color_data = 12'b111011101110;
20'b01000110000100011110: color_data = 12'b111111111111;
20'b01000110000100011111: color_data = 12'b111011101110;
20'b01000110000100100000: color_data = 12'b111011101110;
20'b01000110000100100010: color_data = 12'b111011101110;
20'b01000110000100100011: color_data = 12'b111011101110;
20'b01000110000100100100: color_data = 12'b111011101110;
20'b01000110000100100101: color_data = 12'b111011101110;
20'b01000110000100100110: color_data = 12'b111111111111;
20'b01000110000100101101: color_data = 12'b111011101110;
20'b01000110000100101110: color_data = 12'b111111111111;
20'b01000110000100101111: color_data = 12'b111011101110;
20'b01000110000100110000: color_data = 12'b111011101110;
20'b01000110000100110010: color_data = 12'b111011101110;
20'b01000110000100110011: color_data = 12'b111011101110;
20'b01000110000100110100: color_data = 12'b111011101110;
20'b01000110000100110101: color_data = 12'b111011101110;
20'b01000110000100110110: color_data = 12'b111111111111;
20'b01000110000100111000: color_data = 12'b111011101110;
20'b01000110000100111001: color_data = 12'b111111111111;
20'b01000110000100111010: color_data = 12'b111011101110;
20'b01000110000100111011: color_data = 12'b111011101110;
20'b01000110000100111100: color_data = 12'b111111111111;
20'b01000110000101000010: color_data = 12'b111011101110;
20'b01000110000101000011: color_data = 12'b111011101110;
20'b01000110000101000100: color_data = 12'b111011101110;
20'b01000110000101000101: color_data = 12'b111011101110;
20'b01000110000101000110: color_data = 12'b111011101110;
20'b01000110000101001000: color_data = 12'b111011101110;
20'b01000110000101001001: color_data = 12'b111011101110;
20'b01000110000101001010: color_data = 12'b111011101110;
20'b01000110000101001011: color_data = 12'b111011101110;
20'b01000110000101001100: color_data = 12'b111011101110;
20'b01000110000101101110: color_data = 12'b111011101110;
20'b01000110000101101111: color_data = 12'b111011101110;
20'b01000110000101110000: color_data = 12'b111011101110;
20'b01000110000101110001: color_data = 12'b111111111111;
20'b01000110000101110010: color_data = 12'b111011101110;
20'b01000110000101110100: color_data = 12'b111011101110;
20'b01000110000101110101: color_data = 12'b111011101110;
20'b01000110000101110110: color_data = 12'b111011101110;
20'b01000110000101110111: color_data = 12'b111011101110;
20'b01000110000101111000: color_data = 12'b111011101110;
20'b01000110000101111111: color_data = 12'b111011101110;
20'b01000110000110000000: color_data = 12'b111011101110;
20'b01000110000110000001: color_data = 12'b111011101110;
20'b01000110000110000010: color_data = 12'b111011101110;
20'b01000110000110000100: color_data = 12'b111011101110;
20'b01000110000110000101: color_data = 12'b111011101110;
20'b01000110000110000110: color_data = 12'b111011101110;
20'b01000110000110000111: color_data = 12'b111011101110;
20'b01000110000110001000: color_data = 12'b111011101110;
20'b01000110010011101011: color_data = 12'b111011101110;
20'b01000110010011101100: color_data = 12'b111011101110;
20'b01000110010011101101: color_data = 12'b111011101110;
20'b01000110010011101110: color_data = 12'b111111111111;
20'b01000110010011101111: color_data = 12'b111011101110;
20'b01000110010011110001: color_data = 12'b111011101110;
20'b01000110010011110010: color_data = 12'b111011101110;
20'b01000110010011110011: color_data = 12'b111011101110;
20'b01000110010011110100: color_data = 12'b111111111111;
20'b01000110010011110101: color_data = 12'b111011101110;
20'b01000110010100000111: color_data = 12'b111011101110;
20'b01000110010100001000: color_data = 12'b111011101110;
20'b01000110010100001001: color_data = 12'b111011101110;
20'b01000110010100001010: color_data = 12'b111011101110;
20'b01000110010100001011: color_data = 12'b111011101110;
20'b01000110010100001101: color_data = 12'b111011101110;
20'b01000110010100001110: color_data = 12'b111011101110;
20'b01000110010100001111: color_data = 12'b111011101110;
20'b01000110010100010000: color_data = 12'b111011101110;
20'b01000110010100010111: color_data = 12'b111011101110;
20'b01000110010100011000: color_data = 12'b111011101110;
20'b01000110010100011001: color_data = 12'b111011101110;
20'b01000110010100011010: color_data = 12'b111011101110;
20'b01000110010100011011: color_data = 12'b111011101110;
20'b01000110010100011101: color_data = 12'b111011101110;
20'b01000110010100011110: color_data = 12'b111011101110;
20'b01000110010100011111: color_data = 12'b111111111111;
20'b01000110010100100000: color_data = 12'b111011101110;
20'b01000110010100100010: color_data = 12'b111111111111;
20'b01000110010100100011: color_data = 12'b111011101110;
20'b01000110010100100100: color_data = 12'b111011101110;
20'b01000110010100100101: color_data = 12'b111111111111;
20'b01000110010100100110: color_data = 12'b111011101110;
20'b01000110010100101101: color_data = 12'b111011101110;
20'b01000110010100101110: color_data = 12'b111011101110;
20'b01000110010100101111: color_data = 12'b111111111111;
20'b01000110010100110000: color_data = 12'b111011101110;
20'b01000110010100110010: color_data = 12'b111111111111;
20'b01000110010100110011: color_data = 12'b111011101110;
20'b01000110010100110100: color_data = 12'b111011101110;
20'b01000110010100110101: color_data = 12'b111111111111;
20'b01000110010100110110: color_data = 12'b111011101110;
20'b01000110010100111000: color_data = 12'b111111111111;
20'b01000110010100111001: color_data = 12'b111011101110;
20'b01000110010100111010: color_data = 12'b111011101110;
20'b01000110010100111011: color_data = 12'b111011101110;
20'b01000110010100111100: color_data = 12'b111011101110;
20'b01000110010101000010: color_data = 12'b111011101110;
20'b01000110010101000011: color_data = 12'b111011101110;
20'b01000110010101000100: color_data = 12'b111011101110;
20'b01000110010101000101: color_data = 12'b111011101110;
20'b01000110010101000110: color_data = 12'b111011101110;
20'b01000110010101001000: color_data = 12'b111011101110;
20'b01000110010101001001: color_data = 12'b111011101110;
20'b01000110010101001010: color_data = 12'b111011101110;
20'b01000110010101001011: color_data = 12'b111011101110;
20'b01000110010101001100: color_data = 12'b111011101110;
20'b01000110010101101110: color_data = 12'b111111111111;
20'b01000110010101101111: color_data = 12'b111011101110;
20'b01000110010101110000: color_data = 12'b111111111111;
20'b01000110010101110001: color_data = 12'b111011101110;
20'b01000110010101110010: color_data = 12'b111111111111;
20'b01000110010101110100: color_data = 12'b111011101110;
20'b01000110010101110101: color_data = 12'b111011101110;
20'b01000110010101110110: color_data = 12'b111011101110;
20'b01000110010101110111: color_data = 12'b111011101110;
20'b01000110010101111000: color_data = 12'b111011101110;
20'b01000110010101111111: color_data = 12'b111011101110;
20'b01000110010110000000: color_data = 12'b111011101110;
20'b01000110010110000001: color_data = 12'b111111111111;
20'b01000110010110000010: color_data = 12'b111011101110;
20'b01000110010110000100: color_data = 12'b111011101110;
20'b01000110010110000101: color_data = 12'b111011101110;
20'b01000110010110000110: color_data = 12'b111111111111;
20'b01000110010110000111: color_data = 12'b111011101110;
20'b01000110010110001000: color_data = 12'b111111111111;
20'b01000110100011101011: color_data = 12'b111011101110;
20'b01000110100011101100: color_data = 12'b111111111111;
20'b01000110100011101101: color_data = 12'b111011101110;
20'b01000110100011101110: color_data = 12'b111011101110;
20'b01000110100011101111: color_data = 12'b111111111111;
20'b01000110100011110001: color_data = 12'b111011101110;
20'b01000110100011110010: color_data = 12'b111011101110;
20'b01000110100011110011: color_data = 12'b111011101110;
20'b01000110100011110100: color_data = 12'b111011101110;
20'b01000110100011110101: color_data = 12'b111011101110;
20'b01000110100100000111: color_data = 12'b111011101110;
20'b01000110100100001000: color_data = 12'b111011101110;
20'b01000110100100001001: color_data = 12'b111011101110;
20'b01000110100100001010: color_data = 12'b111011101110;
20'b01000110100100001011: color_data = 12'b111111111111;
20'b01000110100100001101: color_data = 12'b111011101110;
20'b01000110100100001110: color_data = 12'b111111111111;
20'b01000110100100001111: color_data = 12'b111011101110;
20'b01000110100100010000: color_data = 12'b111011101110;
20'b01000110100100010111: color_data = 12'b111111111111;
20'b01000110100100011000: color_data = 12'b111011101110;
20'b01000110100100011001: color_data = 12'b111011101110;
20'b01000110100100011010: color_data = 12'b111011101110;
20'b01000110100100011011: color_data = 12'b111011101110;
20'b01000110100100011101: color_data = 12'b111011101110;
20'b01000110100100011110: color_data = 12'b111011101110;
20'b01000110100100011111: color_data = 12'b111011101110;
20'b01000110100100100000: color_data = 12'b111011101110;
20'b01000110100100100010: color_data = 12'b111011101110;
20'b01000110100100100011: color_data = 12'b111111111111;
20'b01000110100100100100: color_data = 12'b111011101110;
20'b01000110100100100101: color_data = 12'b111011101110;
20'b01000110100100100110: color_data = 12'b111011101110;
20'b01000110100100101101: color_data = 12'b111011101110;
20'b01000110100100101110: color_data = 12'b111011101110;
20'b01000110100100101111: color_data = 12'b111011101110;
20'b01000110100100110000: color_data = 12'b111011101110;
20'b01000110100100110010: color_data = 12'b111011101110;
20'b01000110100100110011: color_data = 12'b111111111111;
20'b01000110100100110100: color_data = 12'b111011101110;
20'b01000110100100110101: color_data = 12'b111011101110;
20'b01000110100100110110: color_data = 12'b111011101110;
20'b01000110100100111000: color_data = 12'b111011101110;
20'b01000110100100111001: color_data = 12'b111011101110;
20'b01000110100100111010: color_data = 12'b111011101110;
20'b01000110100100111011: color_data = 12'b111111111111;
20'b01000110100100111100: color_data = 12'b111011101110;
20'b01000110100101000010: color_data = 12'b111011101110;
20'b01000110100101000011: color_data = 12'b111011101110;
20'b01000110100101000100: color_data = 12'b111011101110;
20'b01000110100101000101: color_data = 12'b111011101110;
20'b01000110100101000110: color_data = 12'b111011101110;
20'b01000110100101001000: color_data = 12'b111011101110;
20'b01000110100101001001: color_data = 12'b111011101110;
20'b01000110100101001010: color_data = 12'b111011101110;
20'b01000110100101001011: color_data = 12'b111011101110;
20'b01000110100101001100: color_data = 12'b111011101110;
20'b01000110100101101110: color_data = 12'b111011101110;
20'b01000110100101101111: color_data = 12'b111011101110;
20'b01000110100101110000: color_data = 12'b111011101110;
20'b01000110100101110001: color_data = 12'b111011101110;
20'b01000110100101110010: color_data = 12'b111011101110;
20'b01000110100101110100: color_data = 12'b111111111111;
20'b01000110100101110101: color_data = 12'b111011101110;
20'b01000110100101110110: color_data = 12'b111011101110;
20'b01000110100101110111: color_data = 12'b111011101110;
20'b01000110100101111000: color_data = 12'b111011101110;
20'b01000110100101111111: color_data = 12'b111111111111;
20'b01000110100110000000: color_data = 12'b111111111111;
20'b01000110100110000001: color_data = 12'b111011101110;
20'b01000110100110000010: color_data = 12'b111111111111;
20'b01000110100110000100: color_data = 12'b111011101110;
20'b01000110100110000101: color_data = 12'b111011101110;
20'b01000110100110000110: color_data = 12'b111011101110;
20'b01000110100110000111: color_data = 12'b111011101110;
20'b01000110100110001000: color_data = 12'b111011101110;
20'b01000110110011101011: color_data = 12'b111011101110;
20'b01000110110011101100: color_data = 12'b111011101110;
20'b01000110110011101101: color_data = 12'b111011101110;
20'b01000110110011101110: color_data = 12'b111011101110;
20'b01000110110011101111: color_data = 12'b111011101110;
20'b01000110110011110001: color_data = 12'b111011101110;
20'b01000110110011110010: color_data = 12'b111011101110;
20'b01000110110011110011: color_data = 12'b111011101110;
20'b01000110110011110100: color_data = 12'b111111111111;
20'b01000110110011110101: color_data = 12'b111011101110;
20'b01000110110100000111: color_data = 12'b111011101110;
20'b01000110110100001000: color_data = 12'b111011101110;
20'b01000110110100001001: color_data = 12'b111011101110;
20'b01000110110100001010: color_data = 12'b111011101110;
20'b01000110110100001011: color_data = 12'b111011101110;
20'b01000110110100001101: color_data = 12'b111011101110;
20'b01000110110100001110: color_data = 12'b111011101110;
20'b01000110110100001111: color_data = 12'b111011101110;
20'b01000110110100010000: color_data = 12'b111011101110;
20'b01000110110100010111: color_data = 12'b111011101110;
20'b01000110110100011000: color_data = 12'b111011101110;
20'b01000110110100011001: color_data = 12'b111011101110;
20'b01000110110100011010: color_data = 12'b111011101110;
20'b01000110110100011011: color_data = 12'b111011101110;
20'b01000110110100011101: color_data = 12'b111011101110;
20'b01000110110100011110: color_data = 12'b111011101110;
20'b01000110110100011111: color_data = 12'b111011101110;
20'b01000110110100100000: color_data = 12'b111011101110;
20'b01000110110100100010: color_data = 12'b111011101110;
20'b01000110110100100011: color_data = 12'b111011101110;
20'b01000110110100100100: color_data = 12'b111111111111;
20'b01000110110100100101: color_data = 12'b111011101110;
20'b01000110110100100110: color_data = 12'b111011101110;
20'b01000110110100101101: color_data = 12'b111011101110;
20'b01000110110100101110: color_data = 12'b111011101110;
20'b01000110110100101111: color_data = 12'b111011101110;
20'b01000110110100110000: color_data = 12'b111011101110;
20'b01000110110100110010: color_data = 12'b111011101110;
20'b01000110110100110011: color_data = 12'b111011101110;
20'b01000110110100110100: color_data = 12'b111111111111;
20'b01000110110100110101: color_data = 12'b111011101110;
20'b01000110110100110110: color_data = 12'b111011101110;
20'b01000110110100111000: color_data = 12'b111011101110;
20'b01000110110100111001: color_data = 12'b111011101110;
20'b01000110110100111010: color_data = 12'b111111111111;
20'b01000110110100111011: color_data = 12'b111011101110;
20'b01000110110100111100: color_data = 12'b111011101110;
20'b01000110110101000010: color_data = 12'b111011101110;
20'b01000110110101000011: color_data = 12'b111111111111;
20'b01000110110101000100: color_data = 12'b111011101110;
20'b01000110110101000101: color_data = 12'b111011101110;
20'b01000110110101000110: color_data = 12'b111011101110;
20'b01000110110101001000: color_data = 12'b111011101110;
20'b01000110110101001001: color_data = 12'b111011101110;
20'b01000110110101001010: color_data = 12'b111011101110;
20'b01000110110101001011: color_data = 12'b111011101110;
20'b01000110110101001100: color_data = 12'b111111111111;
20'b01000110110101101110: color_data = 12'b111011101110;
20'b01000110110101101111: color_data = 12'b111011101110;
20'b01000110110101110000: color_data = 12'b111011101110;
20'b01000110110101110001: color_data = 12'b111011101110;
20'b01000110110101110010: color_data = 12'b111111111111;
20'b01000110110101110100: color_data = 12'b111011101110;
20'b01000110110101110101: color_data = 12'b111011101110;
20'b01000110110101110110: color_data = 12'b111011101110;
20'b01000110110101110111: color_data = 12'b111011101110;
20'b01000110110101111000: color_data = 12'b111011101110;
20'b01000110110101111111: color_data = 12'b111011101110;
20'b01000110110110000000: color_data = 12'b111011101110;
20'b01000110110110000001: color_data = 12'b111011101110;
20'b01000110110110000010: color_data = 12'b111011101110;
20'b01000110110110000100: color_data = 12'b111111111111;
20'b01000110110110000101: color_data = 12'b111011101110;
20'b01000110110110000110: color_data = 12'b111011101110;
20'b01000110110110000111: color_data = 12'b111011101110;
20'b01000110110110001000: color_data = 12'b111011101110;
20'b01000111000011101011: color_data = 12'b111011101110;
20'b01000111000011101100: color_data = 12'b111111111111;
20'b01000111000011101101: color_data = 12'b111011101110;
20'b01000111000011101110: color_data = 12'b111011101110;
20'b01000111000011101111: color_data = 12'b111111111111;
20'b01000111000011110001: color_data = 12'b111011101110;
20'b01000111000011110010: color_data = 12'b111111111111;
20'b01000111000011110011: color_data = 12'b111011101110;
20'b01000111000011110100: color_data = 12'b111011101110;
20'b01000111000011110101: color_data = 12'b111011101110;
20'b01000111000100000111: color_data = 12'b111011101110;
20'b01000111000100001000: color_data = 12'b111011101110;
20'b01000111000100001001: color_data = 12'b111111111111;
20'b01000111000100001010: color_data = 12'b111011101110;
20'b01000111000100001011: color_data = 12'b111011101110;
20'b01000111000100001101: color_data = 12'b111011101110;
20'b01000111000100001110: color_data = 12'b111011101110;
20'b01000111000100001111: color_data = 12'b111011101110;
20'b01000111000100010000: color_data = 12'b111011101110;
20'b01000111000100010111: color_data = 12'b111011101110;
20'b01000111000100011000: color_data = 12'b111011101110;
20'b01000111000100011001: color_data = 12'b111011101110;
20'b01000111000100011010: color_data = 12'b111111111111;
20'b01000111000100011011: color_data = 12'b111011101110;
20'b01000111000100011101: color_data = 12'b111011101110;
20'b01000111000100011110: color_data = 12'b111011101110;
20'b01000111000100011111: color_data = 12'b111011101110;
20'b01000111000100100000: color_data = 12'b111011101110;
20'b01000111000100100010: color_data = 12'b111011101110;
20'b01000111000100100011: color_data = 12'b111011101110;
20'b01000111000100100100: color_data = 12'b111011101110;
20'b01000111000100100101: color_data = 12'b111011101110;
20'b01000111000100100110: color_data = 12'b111011101110;
20'b01000111000100101101: color_data = 12'b111011101110;
20'b01000111000100101110: color_data = 12'b111111111111;
20'b01000111000100101111: color_data = 12'b111011101110;
20'b01000111000100110000: color_data = 12'b111011101110;
20'b01000111000100110010: color_data = 12'b111011101110;
20'b01000111000100110011: color_data = 12'b111011101110;
20'b01000111000100110100: color_data = 12'b111011101110;
20'b01000111000100110101: color_data = 12'b111011101110;
20'b01000111000100110110: color_data = 12'b111011101110;
20'b01000111000100111000: color_data = 12'b111011101110;
20'b01000111000100111001: color_data = 12'b111011101110;
20'b01000111000100111010: color_data = 12'b111011101110;
20'b01000111000100111011: color_data = 12'b111011101110;
20'b01000111000100111100: color_data = 12'b111011101110;
20'b01000111000101000010: color_data = 12'b111011101110;
20'b01000111000101000011: color_data = 12'b111011101110;
20'b01000111000101000100: color_data = 12'b111111111111;
20'b01000111000101000101: color_data = 12'b111011101110;
20'b01000111000101000110: color_data = 12'b111111111111;
20'b01000111000101001000: color_data = 12'b111011101110;
20'b01000111000101001001: color_data = 12'b111011101110;
20'b01000111000101001010: color_data = 12'b111011101110;
20'b01000111000101001011: color_data = 12'b111011101110;
20'b01000111000101001100: color_data = 12'b111011101110;
20'b01000111000101101110: color_data = 12'b111111111111;
20'b01000111000101101111: color_data = 12'b111011101110;
20'b01000111000101110000: color_data = 12'b111011101110;
20'b01000111000101110001: color_data = 12'b111011101110;
20'b01000111000101110010: color_data = 12'b111011101110;
20'b01000111000101110100: color_data = 12'b111011101110;
20'b01000111000101110101: color_data = 12'b111011101110;
20'b01000111000101110110: color_data = 12'b111011101110;
20'b01000111000101110111: color_data = 12'b111011101110;
20'b01000111000101111000: color_data = 12'b111011101110;
20'b01000111000101111111: color_data = 12'b111011101110;
20'b01000111000110000000: color_data = 12'b111011101110;
20'b01000111000110000001: color_data = 12'b111011101110;
20'b01000111000110000010: color_data = 12'b111011101110;
20'b01000111000110000100: color_data = 12'b111011101110;
20'b01000111000110000101: color_data = 12'b111011101110;
20'b01000111000110000110: color_data = 12'b111011101110;
20'b01000111000110000111: color_data = 12'b111011101110;
20'b01000111000110001000: color_data = 12'b111011101110;
20'b01000111100011110001: color_data = 12'b111111111111;
20'b01000111100011110010: color_data = 12'b111011101110;
20'b01000111100011110011: color_data = 12'b111111111111;
20'b01000111100011110100: color_data = 12'b111011101110;
20'b01000111100011110101: color_data = 12'b111011101110;
20'b01000111100011110111: color_data = 12'b111011101110;
20'b01000111100011111000: color_data = 12'b111011101110;
20'b01000111100011111001: color_data = 12'b111011101110;
20'b01000111100011111010: color_data = 12'b111111111111;
20'b01000111100011111100: color_data = 12'b111011101110;
20'b01000111100011111101: color_data = 12'b111011101110;
20'b01000111100011111110: color_data = 12'b111011101110;
20'b01000111100011111111: color_data = 12'b111011101110;
20'b01000111100100000000: color_data = 12'b111011101110;
20'b01000111100100000010: color_data = 12'b111111111111;
20'b01000111100100000011: color_data = 12'b111011101110;
20'b01000111100100000100: color_data = 12'b111011101110;
20'b01000111100100000101: color_data = 12'b111011101110;
20'b01000111100100000111: color_data = 12'b111011101110;
20'b01000111100100001000: color_data = 12'b111011101110;
20'b01000111100100001001: color_data = 12'b111011101110;
20'b01000111100100001010: color_data = 12'b111011101110;
20'b01000111100100001011: color_data = 12'b111111111111;
20'b01000111100100011101: color_data = 12'b111011101110;
20'b01000111100100011110: color_data = 12'b111011101110;
20'b01000111100100011111: color_data = 12'b111011101110;
20'b01000111100100100000: color_data = 12'b111011101110;
20'b01000111100100100010: color_data = 12'b111011101110;
20'b01000111100100100011: color_data = 12'b111011101110;
20'b01000111100100100100: color_data = 12'b111011101110;
20'b01000111100100100101: color_data = 12'b111011101110;
20'b01000111100100100110: color_data = 12'b111011101110;
20'b01000111100100101000: color_data = 12'b111011101110;
20'b01000111100100101001: color_data = 12'b111011101110;
20'b01000111100100101010: color_data = 12'b111011101110;
20'b01000111100100101011: color_data = 12'b111011101110;
20'b01000111100100101101: color_data = 12'b111011101110;
20'b01000111100100101110: color_data = 12'b111011101110;
20'b01000111100100101111: color_data = 12'b111011101110;
20'b01000111100100110000: color_data = 12'b111011101110;
20'b01000111100100110010: color_data = 12'b111011101110;
20'b01000111100100110011: color_data = 12'b111011101110;
20'b01000111100100110100: color_data = 12'b111011101110;
20'b01000111100100110101: color_data = 12'b111011101110;
20'b01000111100100110110: color_data = 12'b111011101110;
20'b01000111100101000010: color_data = 12'b111011101110;
20'b01000111100101000011: color_data = 12'b111011101110;
20'b01000111100101000100: color_data = 12'b111011101110;
20'b01000111100101000101: color_data = 12'b111011101110;
20'b01000111100101000110: color_data = 12'b111111111111;
20'b01000111100101001000: color_data = 12'b111011101110;
20'b01000111100101001001: color_data = 12'b111011101110;
20'b01000111100101001010: color_data = 12'b111011101110;
20'b01000111100101001011: color_data = 12'b111011101110;
20'b01000111100101001100: color_data = 12'b111011101110;
20'b01000111100101001110: color_data = 12'b111011101110;
20'b01000111100101001111: color_data = 12'b111011101110;
20'b01000111100101010000: color_data = 12'b111011101110;
20'b01000111100101010001: color_data = 12'b111011101110;
20'b01000111100101010011: color_data = 12'b111011101110;
20'b01000111100101010100: color_data = 12'b111011101110;
20'b01000111100101010101: color_data = 12'b111011101110;
20'b01000111100101010110: color_data = 12'b111111111111;
20'b01000111100101011000: color_data = 12'b111011101110;
20'b01000111100101011001: color_data = 12'b111111111111;
20'b01000111100101011010: color_data = 12'b111011101110;
20'b01000111100101011011: color_data = 12'b111011101110;
20'b01000111100101011100: color_data = 12'b111011101110;
20'b01000111100101011110: color_data = 12'b111011101110;
20'b01000111100101011111: color_data = 12'b111011101110;
20'b01000111100101100000: color_data = 12'b111011101110;
20'b01000111100101100001: color_data = 12'b111011101110;
20'b01000111100101100011: color_data = 12'b111011101110;
20'b01000111100101100100: color_data = 12'b111011101110;
20'b01000111100101100101: color_data = 12'b111011101110;
20'b01000111100101100110: color_data = 12'b111111111111;
20'b01000111100101100111: color_data = 12'b111011101110;
20'b01000111100101101110: color_data = 12'b111011101110;
20'b01000111100101101111: color_data = 12'b111011101110;
20'b01000111100101110000: color_data = 12'b111011101110;
20'b01000111100101110001: color_data = 12'b111011101110;
20'b01000111100101110010: color_data = 12'b111011101110;
20'b01000111100101110100: color_data = 12'b111011101110;
20'b01000111100101110101: color_data = 12'b111011101110;
20'b01000111100101110110: color_data = 12'b111011101110;
20'b01000111100101110111: color_data = 12'b111011101110;
20'b01000111100101111000: color_data = 12'b111011101110;
20'b01000111100110000100: color_data = 12'b111011101110;
20'b01000111100110000101: color_data = 12'b111011101110;
20'b01000111100110000110: color_data = 12'b111011101110;
20'b01000111100110000111: color_data = 12'b111011101110;
20'b01000111100110001000: color_data = 12'b111011101110;
20'b01000111100110001010: color_data = 12'b111011101110;
20'b01000111100110001011: color_data = 12'b111011101110;
20'b01000111100110001100: color_data = 12'b111011101110;
20'b01000111100110001101: color_data = 12'b111011101110;
20'b01000111100110001110: color_data = 12'b111111111111;
20'b01000111110011110001: color_data = 12'b111011101110;
20'b01000111110011110010: color_data = 12'b111011101110;
20'b01000111110011110011: color_data = 12'b111011101110;
20'b01000111110011110100: color_data = 12'b111011101110;
20'b01000111110011110101: color_data = 12'b111011101110;
20'b01000111110011110111: color_data = 12'b111011101110;
20'b01000111110011111000: color_data = 12'b111011101110;
20'b01000111110011111001: color_data = 12'b111111111111;
20'b01000111110011111010: color_data = 12'b111011101110;
20'b01000111110011111100: color_data = 12'b111011101110;
20'b01000111110011111101: color_data = 12'b111011101110;
20'b01000111110011111110: color_data = 12'b111011101110;
20'b01000111110011111111: color_data = 12'b111011101110;
20'b01000111110100000000: color_data = 12'b111011101110;
20'b01000111110100000010: color_data = 12'b111011101110;
20'b01000111110100000011: color_data = 12'b111011101110;
20'b01000111110100000100: color_data = 12'b111011101110;
20'b01000111110100000101: color_data = 12'b111011101110;
20'b01000111110100000111: color_data = 12'b111011101110;
20'b01000111110100001000: color_data = 12'b111011101110;
20'b01000111110100001001: color_data = 12'b111011101110;
20'b01000111110100001010: color_data = 12'b111011101110;
20'b01000111110100001011: color_data = 12'b111011101110;
20'b01000111110100011101: color_data = 12'b111011101110;
20'b01000111110100011110: color_data = 12'b111011101110;
20'b01000111110100011111: color_data = 12'b111011101110;
20'b01000111110100100000: color_data = 12'b111011101110;
20'b01000111110100100010: color_data = 12'b111011101110;
20'b01000111110100100011: color_data = 12'b111011101110;
20'b01000111110100100100: color_data = 12'b111011101110;
20'b01000111110100100101: color_data = 12'b111011101110;
20'b01000111110100100110: color_data = 12'b111011101110;
20'b01000111110100101000: color_data = 12'b111011101110;
20'b01000111110100101001: color_data = 12'b111011101110;
20'b01000111110100101010: color_data = 12'b111011101110;
20'b01000111110100101011: color_data = 12'b111011101110;
20'b01000111110100101101: color_data = 12'b111111111111;
20'b01000111110100101110: color_data = 12'b111011101110;
20'b01000111110100101111: color_data = 12'b111011101110;
20'b01000111110100110000: color_data = 12'b111011101110;
20'b01000111110100110010: color_data = 12'b111011101110;
20'b01000111110100110011: color_data = 12'b111011101110;
20'b01000111110100110100: color_data = 12'b111011101110;
20'b01000111110100110101: color_data = 12'b111011101110;
20'b01000111110100110110: color_data = 12'b111011101110;
20'b01000111110101000010: color_data = 12'b111011101110;
20'b01000111110101000011: color_data = 12'b111011101110;
20'b01000111110101000100: color_data = 12'b111011101110;
20'b01000111110101000101: color_data = 12'b111011101110;
20'b01000111110101000110: color_data = 12'b111011101110;
20'b01000111110101001000: color_data = 12'b111011101110;
20'b01000111110101001001: color_data = 12'b111011101110;
20'b01000111110101001010: color_data = 12'b111011101110;
20'b01000111110101001011: color_data = 12'b111011101110;
20'b01000111110101001100: color_data = 12'b111011101110;
20'b01000111110101001110: color_data = 12'b111011101110;
20'b01000111110101001111: color_data = 12'b111011101110;
20'b01000111110101010000: color_data = 12'b111011101110;
20'b01000111110101010001: color_data = 12'b111011101110;
20'b01000111110101010011: color_data = 12'b111011101110;
20'b01000111110101010100: color_data = 12'b111011101110;
20'b01000111110101010101: color_data = 12'b111011101110;
20'b01000111110101010110: color_data = 12'b111011101110;
20'b01000111110101011000: color_data = 12'b111011101110;
20'b01000111110101011001: color_data = 12'b111011101110;
20'b01000111110101011010: color_data = 12'b111011101110;
20'b01000111110101011011: color_data = 12'b111011101110;
20'b01000111110101011100: color_data = 12'b111011101110;
20'b01000111110101011110: color_data = 12'b111011101110;
20'b01000111110101011111: color_data = 12'b111011101110;
20'b01000111110101100000: color_data = 12'b111011101110;
20'b01000111110101100001: color_data = 12'b111011101110;
20'b01000111110101100011: color_data = 12'b111011101110;
20'b01000111110101100100: color_data = 12'b111011101110;
20'b01000111110101100101: color_data = 12'b111011101110;
20'b01000111110101100110: color_data = 12'b111011101110;
20'b01000111110101100111: color_data = 12'b111011101110;
20'b01000111110101101110: color_data = 12'b111011101110;
20'b01000111110101101111: color_data = 12'b111011101110;
20'b01000111110101110000: color_data = 12'b111011101110;
20'b01000111110101110001: color_data = 12'b111011101110;
20'b01000111110101110010: color_data = 12'b111011101110;
20'b01000111110101110100: color_data = 12'b111011101110;
20'b01000111110101110101: color_data = 12'b111111111111;
20'b01000111110101110110: color_data = 12'b111011101110;
20'b01000111110101110111: color_data = 12'b111011101110;
20'b01000111110101111000: color_data = 12'b111011101110;
20'b01000111110110000100: color_data = 12'b111011101110;
20'b01000111110110000101: color_data = 12'b111111111111;
20'b01000111110110000110: color_data = 12'b111011101110;
20'b01000111110110000111: color_data = 12'b111011101110;
20'b01000111110110001000: color_data = 12'b111011101110;
20'b01000111110110001010: color_data = 12'b111011101110;
20'b01000111110110001011: color_data = 12'b111011101110;
20'b01000111110110001100: color_data = 12'b111011101110;
20'b01000111110110001101: color_data = 12'b111011101110;
20'b01000111110110001110: color_data = 12'b111011101110;
20'b01001000000011110001: color_data = 12'b111011101110;
20'b01001000000011110010: color_data = 12'b111011101110;
20'b01001000000011110011: color_data = 12'b111011101110;
20'b01001000000011110100: color_data = 12'b111011101110;
20'b01001000000011110101: color_data = 12'b111011101110;
20'b01001000000011110111: color_data = 12'b111011101110;
20'b01001000000011111000: color_data = 12'b111111111111;
20'b01001000000011111001: color_data = 12'b111011101110;
20'b01001000000011111010: color_data = 12'b111011101110;
20'b01001000000011111100: color_data = 12'b111011101110;
20'b01001000000011111101: color_data = 12'b111011101110;
20'b01001000000011111110: color_data = 12'b111011101110;
20'b01001000000011111111: color_data = 12'b111011101110;
20'b01001000000100000000: color_data = 12'b111011101110;
20'b01001000000100000010: color_data = 12'b111011101110;
20'b01001000000100000011: color_data = 12'b111011101110;
20'b01001000000100000100: color_data = 12'b111011101110;
20'b01001000000100000101: color_data = 12'b111011101110;
20'b01001000000100000111: color_data = 12'b111011101110;
20'b01001000000100001000: color_data = 12'b111011101110;
20'b01001000000100001001: color_data = 12'b111011101110;
20'b01001000000100001010: color_data = 12'b111011101110;
20'b01001000000100001011: color_data = 12'b111011101110;
20'b01001000000100011101: color_data = 12'b111011101110;
20'b01001000000100011110: color_data = 12'b111011101110;
20'b01001000000100011111: color_data = 12'b111011101110;
20'b01001000000100100000: color_data = 12'b111011101110;
20'b01001000000100100010: color_data = 12'b111011101110;
20'b01001000000100100011: color_data = 12'b111011101110;
20'b01001000000100100100: color_data = 12'b111011101110;
20'b01001000000100100101: color_data = 12'b111111111111;
20'b01001000000100100110: color_data = 12'b111011101110;
20'b01001000000100101000: color_data = 12'b111011101110;
20'b01001000000100101001: color_data = 12'b111011101110;
20'b01001000000100101010: color_data = 12'b111011101110;
20'b01001000000100101011: color_data = 12'b111011101110;
20'b01001000000100101101: color_data = 12'b111011101110;
20'b01001000000100101110: color_data = 12'b111011101110;
20'b01001000000100101111: color_data = 12'b111111111111;
20'b01001000000100110000: color_data = 12'b111011101110;
20'b01001000000100110010: color_data = 12'b111111111111;
20'b01001000000100110011: color_data = 12'b111011101110;
20'b01001000000100110100: color_data = 12'b111011101110;
20'b01001000000100110101: color_data = 12'b111111111111;
20'b01001000000100110110: color_data = 12'b111011101110;
20'b01001000000101000010: color_data = 12'b111011101110;
20'b01001000000101000011: color_data = 12'b111011101110;
20'b01001000000101000100: color_data = 12'b111011101110;
20'b01001000000101000101: color_data = 12'b111011101110;
20'b01001000000101000110: color_data = 12'b111011101110;
20'b01001000000101001000: color_data = 12'b111011101110;
20'b01001000000101001001: color_data = 12'b111011101110;
20'b01001000000101001010: color_data = 12'b111011101110;
20'b01001000000101001011: color_data = 12'b111011101110;
20'b01001000000101001100: color_data = 12'b111011101110;
20'b01001000000101001110: color_data = 12'b111011101110;
20'b01001000000101001111: color_data = 12'b111011101110;
20'b01001000000101010000: color_data = 12'b111111111111;
20'b01001000000101010001: color_data = 12'b111011101110;
20'b01001000000101010011: color_data = 12'b111011101110;
20'b01001000000101010100: color_data = 12'b111011101110;
20'b01001000000101010101: color_data = 12'b111011101110;
20'b01001000000101010110: color_data = 12'b111011101110;
20'b01001000000101011000: color_data = 12'b111011101110;
20'b01001000000101011001: color_data = 12'b111011101110;
20'b01001000000101011010: color_data = 12'b111011101110;
20'b01001000000101011011: color_data = 12'b111011101110;
20'b01001000000101011100: color_data = 12'b111011101110;
20'b01001000000101011110: color_data = 12'b111011101110;
20'b01001000000101011111: color_data = 12'b111011101110;
20'b01001000000101100000: color_data = 12'b111011101110;
20'b01001000000101100001: color_data = 12'b111011101110;
20'b01001000000101100011: color_data = 12'b111011101110;
20'b01001000000101100100: color_data = 12'b111011101110;
20'b01001000000101100101: color_data = 12'b111011101110;
20'b01001000000101100110: color_data = 12'b111011101110;
20'b01001000000101100111: color_data = 12'b111011101110;
20'b01001000000101101110: color_data = 12'b111111111111;
20'b01001000000101101111: color_data = 12'b111011101110;
20'b01001000000101110000: color_data = 12'b111111111111;
20'b01001000000101110001: color_data = 12'b111011101110;
20'b01001000000101110010: color_data = 12'b111011101110;
20'b01001000000101110100: color_data = 12'b111011101110;
20'b01001000000101110101: color_data = 12'b111011101110;
20'b01001000000101110110: color_data = 12'b111011101110;
20'b01001000000101110111: color_data = 12'b111011101110;
20'b01001000000101111000: color_data = 12'b111011101110;
20'b01001000000110000100: color_data = 12'b111011101110;
20'b01001000000110000101: color_data = 12'b111011101110;
20'b01001000000110000110: color_data = 12'b111011101110;
20'b01001000000110000111: color_data = 12'b111011101110;
20'b01001000000110001000: color_data = 12'b111011101110;
20'b01001000000110001010: color_data = 12'b111011101110;
20'b01001000000110001011: color_data = 12'b111011101110;
20'b01001000000110001100: color_data = 12'b111011101110;
20'b01001000000110001101: color_data = 12'b111111111111;
20'b01001000000110001110: color_data = 12'b111011101110;
20'b01001000010011110001: color_data = 12'b111011101110;
20'b01001000010011110010: color_data = 12'b111011101110;
20'b01001000010011110011: color_data = 12'b111111111111;
20'b01001000010011110100: color_data = 12'b111011101110;
20'b01001000010011110101: color_data = 12'b111011101110;
20'b01001000010011110111: color_data = 12'b111011101110;
20'b01001000010011111000: color_data = 12'b111011101110;
20'b01001000010011111001: color_data = 12'b111011101110;
20'b01001000010011111010: color_data = 12'b111111111111;
20'b01001000010011111100: color_data = 12'b111011101110;
20'b01001000010011111101: color_data = 12'b111111111111;
20'b01001000010011111110: color_data = 12'b111011101110;
20'b01001000010011111111: color_data = 12'b111011101110;
20'b01001000010100000000: color_data = 12'b111011101110;
20'b01001000010100000010: color_data = 12'b111011101110;
20'b01001000010100000011: color_data = 12'b111011101110;
20'b01001000010100000100: color_data = 12'b111011101110;
20'b01001000010100000101: color_data = 12'b111011101110;
20'b01001000010100000111: color_data = 12'b111011101110;
20'b01001000010100001000: color_data = 12'b111011101110;
20'b01001000010100001001: color_data = 12'b111011101110;
20'b01001000010100001010: color_data = 12'b111011101110;
20'b01001000010100001011: color_data = 12'b111011101110;
20'b01001000010100011101: color_data = 12'b111011101110;
20'b01001000010100011110: color_data = 12'b111111111111;
20'b01001000010100011111: color_data = 12'b111011101110;
20'b01001000010100100000: color_data = 12'b111011101110;
20'b01001000010100100010: color_data = 12'b111011101110;
20'b01001000010100100011: color_data = 12'b111011101110;
20'b01001000010100100100: color_data = 12'b111111111111;
20'b01001000010100100101: color_data = 12'b111011101110;
20'b01001000010100100110: color_data = 12'b111011101110;
20'b01001000010100101000: color_data = 12'b111011101110;
20'b01001000010100101001: color_data = 12'b111011101110;
20'b01001000010100101010: color_data = 12'b111111111111;
20'b01001000010100101011: color_data = 12'b111011101110;
20'b01001000010100101101: color_data = 12'b111111111111;
20'b01001000010100101110: color_data = 12'b111011101110;
20'b01001000010100101111: color_data = 12'b111011101110;
20'b01001000010100110000: color_data = 12'b111011101110;
20'b01001000010100110010: color_data = 12'b111011101110;
20'b01001000010100110011: color_data = 12'b111011101110;
20'b01001000010100110100: color_data = 12'b111011101110;
20'b01001000010100110101: color_data = 12'b111011101110;
20'b01001000010100110110: color_data = 12'b111011101110;
20'b01001000010101000010: color_data = 12'b111011101110;
20'b01001000010101000011: color_data = 12'b111011101110;
20'b01001000010101000100: color_data = 12'b111011101110;
20'b01001000010101000101: color_data = 12'b111011101110;
20'b01001000010101000110: color_data = 12'b111011101110;
20'b01001000010101001000: color_data = 12'b111111111111;
20'b01001000010101001001: color_data = 12'b111011101110;
20'b01001000010101001010: color_data = 12'b111011101110;
20'b01001000010101001011: color_data = 12'b111011101110;
20'b01001000010101001100: color_data = 12'b111011101110;
20'b01001000010101001110: color_data = 12'b111011101110;
20'b01001000010101001111: color_data = 12'b111011101110;
20'b01001000010101010000: color_data = 12'b111011101110;
20'b01001000010101010001: color_data = 12'b111011101110;
20'b01001000010101010011: color_data = 12'b111111111111;
20'b01001000010101010100: color_data = 12'b111011101110;
20'b01001000010101010101: color_data = 12'b111011101110;
20'b01001000010101010110: color_data = 12'b111011101110;
20'b01001000010101011000: color_data = 12'b111111111111;
20'b01001000010101011001: color_data = 12'b111011101110;
20'b01001000010101011010: color_data = 12'b111011101110;
20'b01001000010101011011: color_data = 12'b111011101110;
20'b01001000010101011100: color_data = 12'b111011101110;
20'b01001000010101011110: color_data = 12'b111011101110;
20'b01001000010101011111: color_data = 12'b111011101110;
20'b01001000010101100000: color_data = 12'b111011101110;
20'b01001000010101100001: color_data = 12'b111011101110;
20'b01001000010101100011: color_data = 12'b111011101110;
20'b01001000010101100100: color_data = 12'b111011101110;
20'b01001000010101100101: color_data = 12'b111011101110;
20'b01001000010101100110: color_data = 12'b111011101110;
20'b01001000010101100111: color_data = 12'b111111111111;
20'b01001000010101101110: color_data = 12'b111011101110;
20'b01001000010101101111: color_data = 12'b111111111111;
20'b01001000010101110000: color_data = 12'b111011101110;
20'b01001000010101110001: color_data = 12'b111011101110;
20'b01001000010101110010: color_data = 12'b111111111111;
20'b01001000010101110100: color_data = 12'b111011101110;
20'b01001000010101110101: color_data = 12'b111111111111;
20'b01001000010101110110: color_data = 12'b111011101110;
20'b01001000010101110111: color_data = 12'b111011101110;
20'b01001000010101111000: color_data = 12'b111011101110;
20'b01001000010110000100: color_data = 12'b111011101110;
20'b01001000010110000101: color_data = 12'b111011101110;
20'b01001000010110000110: color_data = 12'b111011101110;
20'b01001000010110000111: color_data = 12'b111011101110;
20'b01001000010110001000: color_data = 12'b111011101110;
20'b01001000010110001010: color_data = 12'b111011101110;
20'b01001000010110001011: color_data = 12'b111011101110;
20'b01001000010110001100: color_data = 12'b111111111111;
20'b01001000010110001101: color_data = 12'b111011101110;
20'b01001000010110001110: color_data = 12'b111011101110;
20'b01001000100011110001: color_data = 12'b111011101110;
20'b01001000100011110010: color_data = 12'b111011101110;
20'b01001000100011110011: color_data = 12'b111011101110;
20'b01001000100011110100: color_data = 12'b111011101110;
20'b01001000100011110101: color_data = 12'b111011101110;
20'b01001000100011110111: color_data = 12'b111111111111;
20'b01001000100011111000: color_data = 12'b111011101110;
20'b01001000100011111001: color_data = 12'b111011101110;
20'b01001000100011111010: color_data = 12'b111011101110;
20'b01001000100011111100: color_data = 12'b111011101110;
20'b01001000100011111101: color_data = 12'b111011101110;
20'b01001000100011111110: color_data = 12'b111111111111;
20'b01001000100011111111: color_data = 12'b111011101110;
20'b01001000100100000000: color_data = 12'b111011101110;
20'b01001000100100000010: color_data = 12'b111011101110;
20'b01001000100100000011: color_data = 12'b111011101110;
20'b01001000100100000100: color_data = 12'b111011101110;
20'b01001000100100000101: color_data = 12'b111011101110;
20'b01001000100100000111: color_data = 12'b111011101110;
20'b01001000100100001000: color_data = 12'b111011101110;
20'b01001000100100001001: color_data = 12'b111011101110;
20'b01001000100100001010: color_data = 12'b111011101110;
20'b01001000100100001011: color_data = 12'b111011101110;
20'b01001000100100011101: color_data = 12'b111111111111;
20'b01001000100100011110: color_data = 12'b111011101110;
20'b01001000100100011111: color_data = 12'b111011101110;
20'b01001000100100100000: color_data = 12'b111111111111;
20'b01001000100100100010: color_data = 12'b111011101110;
20'b01001000100100100011: color_data = 12'b111111111111;
20'b01001000100100100100: color_data = 12'b111011101110;
20'b01001000100100100101: color_data = 12'b111011101110;
20'b01001000100100100110: color_data = 12'b111111111111;
20'b01001000100100101000: color_data = 12'b111011101110;
20'b01001000100100101001: color_data = 12'b111111111111;
20'b01001000100100101010: color_data = 12'b111011101110;
20'b01001000100100101011: color_data = 12'b111011101110;
20'b01001000100100101101: color_data = 12'b111011101110;
20'b01001000100100101110: color_data = 12'b111011101110;
20'b01001000100100101111: color_data = 12'b111011101110;
20'b01001000100100110000: color_data = 12'b111011101110;
20'b01001000100100110010: color_data = 12'b111011101110;
20'b01001000100100110011: color_data = 12'b111011101110;
20'b01001000100100110100: color_data = 12'b111011101110;
20'b01001000100100110101: color_data = 12'b111011101110;
20'b01001000100100110110: color_data = 12'b111111111111;
20'b01001000100101000010: color_data = 12'b111011101110;
20'b01001000100101000011: color_data = 12'b111011101110;
20'b01001000100101000100: color_data = 12'b111011101110;
20'b01001000100101000101: color_data = 12'b111011101110;
20'b01001000100101000110: color_data = 12'b111011101110;
20'b01001000100101001000: color_data = 12'b111011101110;
20'b01001000100101001001: color_data = 12'b111011101110;
20'b01001000100101001010: color_data = 12'b111111111111;
20'b01001000100101001011: color_data = 12'b111111111111;
20'b01001000100101001100: color_data = 12'b111011101110;
20'b01001000100101001110: color_data = 12'b111011101110;
20'b01001000100101001111: color_data = 12'b111111111111;
20'b01001000100101010000: color_data = 12'b111011101110;
20'b01001000100101010001: color_data = 12'b111111111111;
20'b01001000100101010011: color_data = 12'b111011101110;
20'b01001000100101010100: color_data = 12'b111011101110;
20'b01001000100101010101: color_data = 12'b111011101110;
20'b01001000100101010110: color_data = 12'b111011101110;
20'b01001000100101011000: color_data = 12'b111011101110;
20'b01001000100101011001: color_data = 12'b111011101110;
20'b01001000100101011010: color_data = 12'b111111111111;
20'b01001000100101011011: color_data = 12'b111111111111;
20'b01001000100101011100: color_data = 12'b111011101110;
20'b01001000100101011110: color_data = 12'b111011101110;
20'b01001000100101011111: color_data = 12'b111111111111;
20'b01001000100101100000: color_data = 12'b111111111111;
20'b01001000100101100001: color_data = 12'b111011101110;
20'b01001000100101100011: color_data = 12'b111011101110;
20'b01001000100101100100: color_data = 12'b111111111111;
20'b01001000100101100101: color_data = 12'b111111111111;
20'b01001000100101100110: color_data = 12'b111011101110;
20'b01001000100101100111: color_data = 12'b111011101110;
20'b01001000100101101110: color_data = 12'b111111111111;
20'b01001000100101101111: color_data = 12'b111011101110;
20'b01001000100101110000: color_data = 12'b111011101110;
20'b01001000100101110001: color_data = 12'b111011101110;
20'b01001000100101110010: color_data = 12'b111011101110;
20'b01001000100101110100: color_data = 12'b111011101110;
20'b01001000100101110101: color_data = 12'b111011101110;
20'b01001000100101110110: color_data = 12'b111111111111;
20'b01001000100101110111: color_data = 12'b111011101110;
20'b01001000100101111000: color_data = 12'b111011101110;
20'b01001000100110000100: color_data = 12'b111011101110;
20'b01001000100110000101: color_data = 12'b111011101110;
20'b01001000100110000110: color_data = 12'b111011101110;
20'b01001000100110000111: color_data = 12'b111011101110;
20'b01001000100110001000: color_data = 12'b111111111111;
20'b01001000100110001010: color_data = 12'b111011101110;
20'b01001000100110001011: color_data = 12'b111111111111;
20'b01001000100110001100: color_data = 12'b111011101110;
20'b01001000100110001101: color_data = 12'b111011101110;
20'b01001000100110001110: color_data = 12'b111111111111;
20'b01001001000011110001: color_data = 12'b111011101110;
20'b01001001000011110010: color_data = 12'b111011101110;
20'b01001001000011110011: color_data = 12'b111011101110;
20'b01001001000011110100: color_data = 12'b111011101110;
20'b01001001000011110101: color_data = 12'b111011101110;
20'b01001001000011110111: color_data = 12'b111011101110;
20'b01001001000011111000: color_data = 12'b111011101110;
20'b01001001000011111001: color_data = 12'b111011101110;
20'b01001001000011111010: color_data = 12'b111011101110;
20'b01001001000011111100: color_data = 12'b111011101110;
20'b01001001000011111101: color_data = 12'b111011101110;
20'b01001001000011111110: color_data = 12'b111111111111;
20'b01001001000011111111: color_data = 12'b111011101110;
20'b01001001000100000000: color_data = 12'b111011101110;
20'b01001001000100000010: color_data = 12'b111011101110;
20'b01001001000100000011: color_data = 12'b111011101110;
20'b01001001000100000100: color_data = 12'b111011101110;
20'b01001001000100000101: color_data = 12'b111011101110;
20'b01001001000100000111: color_data = 12'b111011101110;
20'b01001001000100001000: color_data = 12'b111011101110;
20'b01001001000100001001: color_data = 12'b111011101110;
20'b01001001000100001010: color_data = 12'b111011101110;
20'b01001001000100001011: color_data = 12'b111011101110;
20'b01001001000100100010: color_data = 12'b111011101110;
20'b01001001000100100011: color_data = 12'b111111111111;
20'b01001001000100100100: color_data = 12'b111011101110;
20'b01001001000100100101: color_data = 12'b111011101110;
20'b01001001000100100110: color_data = 12'b111011101110;
20'b01001001000100101000: color_data = 12'b111011101110;
20'b01001001000100101001: color_data = 12'b111111111111;
20'b01001001000100101010: color_data = 12'b111011101110;
20'b01001001000100101011: color_data = 12'b111011101110;
20'b01001001000100101101: color_data = 12'b111011101110;
20'b01001001000100101110: color_data = 12'b111011101110;
20'b01001001000100101111: color_data = 12'b111011101110;
20'b01001001000100110000: color_data = 12'b111011101110;
20'b01001001000101000010: color_data = 12'b111011101110;
20'b01001001000101000011: color_data = 12'b111011101110;
20'b01001001000101000100: color_data = 12'b111011101110;
20'b01001001000101000101: color_data = 12'b111011101110;
20'b01001001000101000110: color_data = 12'b111011101110;
20'b01001001000101001000: color_data = 12'b111011101110;
20'b01001001000101001001: color_data = 12'b111011101110;
20'b01001001000101001010: color_data = 12'b111011101110;
20'b01001001000101001011: color_data = 12'b111111111111;
20'b01001001000101001100: color_data = 12'b111011101110;
20'b01001001000101001110: color_data = 12'b111111111111;
20'b01001001000101001111: color_data = 12'b111011101110;
20'b01001001000101010000: color_data = 12'b111011101110;
20'b01001001000101010001: color_data = 12'b111011101110;
20'b01001001000101010011: color_data = 12'b111011101110;
20'b01001001000101010100: color_data = 12'b111011101110;
20'b01001001000101010101: color_data = 12'b111011101110;
20'b01001001000101010110: color_data = 12'b111111111111;
20'b01001001000101011000: color_data = 12'b111011101110;
20'b01001001000101011001: color_data = 12'b111011101110;
20'b01001001000101011010: color_data = 12'b111011101110;
20'b01001001000101011011: color_data = 12'b111111111111;
20'b01001001000101011100: color_data = 12'b111011101110;
20'b01001001000101011110: color_data = 12'b111111111111;
20'b01001001000101011111: color_data = 12'b111011101110;
20'b01001001000101100000: color_data = 12'b111011101110;
20'b01001001000101100001: color_data = 12'b111111111111;
20'b01001001000101100011: color_data = 12'b111011101110;
20'b01001001000101100100: color_data = 12'b111111111111;
20'b01001001000101100101: color_data = 12'b111011101110;
20'b01001001000101100110: color_data = 12'b111011101110;
20'b01001001000101100111: color_data = 12'b111011101110;
20'b01001001000101101110: color_data = 12'b111011101110;
20'b01001001000101101111: color_data = 12'b111011101110;
20'b01001001000101110000: color_data = 12'b111011101110;
20'b01001001000101110001: color_data = 12'b111011101110;
20'b01001001000101110010: color_data = 12'b111011101110;
20'b01001001000101110100: color_data = 12'b111011101110;
20'b01001001000101110101: color_data = 12'b111011101110;
20'b01001001000101110110: color_data = 12'b111111111111;
20'b01001001000101110111: color_data = 12'b111011101110;
20'b01001001000101111000: color_data = 12'b111011101110;
20'b01001001000110001010: color_data = 12'b111011101110;
20'b01001001000110001011: color_data = 12'b111111111111;
20'b01001001000110001100: color_data = 12'b111011101110;
20'b01001001000110001101: color_data = 12'b111011101110;
20'b01001001000110001110: color_data = 12'b111011101110;
20'b01001001000110010000: color_data = 12'b111011101110;
20'b01001001000110010001: color_data = 12'b111011101110;
20'b01001001000110010010: color_data = 12'b111011101110;
20'b01001001000110010011: color_data = 12'b111011101110;
20'b01001001010011110001: color_data = 12'b111111111111;
20'b01001001010011110010: color_data = 12'b111011101110;
20'b01001001010011110011: color_data = 12'b111011101110;
20'b01001001010011110100: color_data = 12'b111011101110;
20'b01001001010011110101: color_data = 12'b111011101110;
20'b01001001010011110111: color_data = 12'b111011101110;
20'b01001001010011111000: color_data = 12'b111011101110;
20'b01001001010011111001: color_data = 12'b111111111111;
20'b01001001010011111010: color_data = 12'b111011101110;
20'b01001001010011111100: color_data = 12'b111011101110;
20'b01001001010011111101: color_data = 12'b111111111111;
20'b01001001010011111110: color_data = 12'b111011101110;
20'b01001001010011111111: color_data = 12'b111011101110;
20'b01001001010100000000: color_data = 12'b111011101110;
20'b01001001010100000010: color_data = 12'b111011101110;
20'b01001001010100000011: color_data = 12'b111011101110;
20'b01001001010100000100: color_data = 12'b111011101110;
20'b01001001010100000101: color_data = 12'b111011101110;
20'b01001001010100000111: color_data = 12'b111011101110;
20'b01001001010100001000: color_data = 12'b111011101110;
20'b01001001010100001001: color_data = 12'b111011101110;
20'b01001001010100001010: color_data = 12'b111011101110;
20'b01001001010100001011: color_data = 12'b111011101110;
20'b01001001010100100010: color_data = 12'b111011101110;
20'b01001001010100100011: color_data = 12'b111011101110;
20'b01001001010100100100: color_data = 12'b111011101110;
20'b01001001010100100101: color_data = 12'b111111111111;
20'b01001001010100100110: color_data = 12'b111011101110;
20'b01001001010100101000: color_data = 12'b111011101110;
20'b01001001010100101001: color_data = 12'b111011101110;
20'b01001001010100101010: color_data = 12'b111111111111;
20'b01001001010100101011: color_data = 12'b111011101110;
20'b01001001010100101101: color_data = 12'b111011101110;
20'b01001001010100101110: color_data = 12'b111111111111;
20'b01001001010100101111: color_data = 12'b111011101110;
20'b01001001010100110000: color_data = 12'b111111111111;
20'b01001001010101000010: color_data = 12'b111011101110;
20'b01001001010101000011: color_data = 12'b111011101110;
20'b01001001010101000100: color_data = 12'b111011101110;
20'b01001001010101000101: color_data = 12'b111011101110;
20'b01001001010101000110: color_data = 12'b111111111111;
20'b01001001010101001000: color_data = 12'b111011101110;
20'b01001001010101001001: color_data = 12'b111011101110;
20'b01001001010101001010: color_data = 12'b111011101110;
20'b01001001010101001011: color_data = 12'b111011101110;
20'b01001001010101001100: color_data = 12'b111011101110;
20'b01001001010101001110: color_data = 12'b111011101110;
20'b01001001010101001111: color_data = 12'b111111111111;
20'b01001001010101010000: color_data = 12'b111011101110;
20'b01001001010101010001: color_data = 12'b111011101110;
20'b01001001010101010011: color_data = 12'b111111111111;
20'b01001001010101010100: color_data = 12'b111011101110;
20'b01001001010101010101: color_data = 12'b111011101110;
20'b01001001010101010110: color_data = 12'b111011101110;
20'b01001001010101011000: color_data = 12'b111011101110;
20'b01001001010101011001: color_data = 12'b111011101110;
20'b01001001010101011010: color_data = 12'b111011101110;
20'b01001001010101011011: color_data = 12'b111011101110;
20'b01001001010101011100: color_data = 12'b111011101110;
20'b01001001010101011110: color_data = 12'b111011101110;
20'b01001001010101011111: color_data = 12'b111111111111;
20'b01001001010101100000: color_data = 12'b111111111111;
20'b01001001010101100001: color_data = 12'b111011101110;
20'b01001001010101100011: color_data = 12'b111011101110;
20'b01001001010101100100: color_data = 12'b111011101110;
20'b01001001010101100101: color_data = 12'b111011101110;
20'b01001001010101100110: color_data = 12'b111011101110;
20'b01001001010101100111: color_data = 12'b111011101110;
20'b01001001010101101110: color_data = 12'b111011101110;
20'b01001001010101101111: color_data = 12'b111011101110;
20'b01001001010101110000: color_data = 12'b111011101110;
20'b01001001010101110001: color_data = 12'b111111111111;
20'b01001001010101110010: color_data = 12'b111011101110;
20'b01001001010101110100: color_data = 12'b111011101110;
20'b01001001010101110101: color_data = 12'b111111111111;
20'b01001001010101110110: color_data = 12'b111011101110;
20'b01001001010101110111: color_data = 12'b111011101110;
20'b01001001010101111000: color_data = 12'b111011101110;
20'b01001001010110001010: color_data = 12'b111011101110;
20'b01001001010110001011: color_data = 12'b111011101110;
20'b01001001010110001100: color_data = 12'b111011101110;
20'b01001001010110001101: color_data = 12'b111111111111;
20'b01001001010110001110: color_data = 12'b111011101110;
20'b01001001010110010000: color_data = 12'b111011101110;
20'b01001001010110010001: color_data = 12'b111011101110;
20'b01001001010110010010: color_data = 12'b111011101110;
20'b01001001010110010011: color_data = 12'b111011101110;
20'b01001001100011110001: color_data = 12'b111011101110;
20'b01001001100011110010: color_data = 12'b111011101110;
20'b01001001100011110011: color_data = 12'b111011101110;
20'b01001001100011110100: color_data = 12'b111011101110;
20'b01001001100011110101: color_data = 12'b111111111111;
20'b01001001100011110111: color_data = 12'b111011101110;
20'b01001001100011111000: color_data = 12'b111011101110;
20'b01001001100011111001: color_data = 12'b111011101110;
20'b01001001100011111010: color_data = 12'b111011101110;
20'b01001001100011111100: color_data = 12'b111111111111;
20'b01001001100011111101: color_data = 12'b111011101110;
20'b01001001100011111110: color_data = 12'b111011101110;
20'b01001001100011111111: color_data = 12'b111011101110;
20'b01001001100100000000: color_data = 12'b111011101110;
20'b01001001100100000010: color_data = 12'b111011101110;
20'b01001001100100000011: color_data = 12'b111011101110;
20'b01001001100100000100: color_data = 12'b111011101110;
20'b01001001100100000101: color_data = 12'b111011101110;
20'b01001001100100000111: color_data = 12'b111011101110;
20'b01001001100100001000: color_data = 12'b111011101110;
20'b01001001100100001001: color_data = 12'b111111111111;
20'b01001001100100001010: color_data = 12'b111011101110;
20'b01001001100100001011: color_data = 12'b111011101110;
20'b01001001100100100010: color_data = 12'b111011101110;
20'b01001001100100100011: color_data = 12'b111011101110;
20'b01001001100100100100: color_data = 12'b111011101110;
20'b01001001100100100101: color_data = 12'b111011101110;
20'b01001001100100100110: color_data = 12'b111011101110;
20'b01001001100100101000: color_data = 12'b111011101110;
20'b01001001100100101001: color_data = 12'b111011101110;
20'b01001001100100101010: color_data = 12'b111011101110;
20'b01001001100100101011: color_data = 12'b111111111111;
20'b01001001100100101101: color_data = 12'b111011101110;
20'b01001001100100101110: color_data = 12'b111011101110;
20'b01001001100100101111: color_data = 12'b111011101110;
20'b01001001100100110000: color_data = 12'b111011101110;
20'b01001001100101000010: color_data = 12'b111011101110;
20'b01001001100101000011: color_data = 12'b111011101110;
20'b01001001100101000100: color_data = 12'b111011101110;
20'b01001001100101000101: color_data = 12'b111111111111;
20'b01001001100101000110: color_data = 12'b111011101110;
20'b01001001100101001000: color_data = 12'b111011101110;
20'b01001001100101001001: color_data = 12'b111011101110;
20'b01001001100101001010: color_data = 12'b111011101110;
20'b01001001100101001011: color_data = 12'b111011101110;
20'b01001001100101001100: color_data = 12'b111011101110;
20'b01001001100101001110: color_data = 12'b111011101110;
20'b01001001100101001111: color_data = 12'b111011101110;
20'b01001001100101010000: color_data = 12'b111011101110;
20'b01001001100101010001: color_data = 12'b111011101110;
20'b01001001100101010011: color_data = 12'b111011101110;
20'b01001001100101010100: color_data = 12'b111011101110;
20'b01001001100101010101: color_data = 12'b111011101110;
20'b01001001100101010110: color_data = 12'b111011101110;
20'b01001001100101011000: color_data = 12'b111011101110;
20'b01001001100101011001: color_data = 12'b111011101110;
20'b01001001100101011010: color_data = 12'b111011101110;
20'b01001001100101011011: color_data = 12'b111011101110;
20'b01001001100101011100: color_data = 12'b111011101110;
20'b01001001100101011110: color_data = 12'b111011101110;
20'b01001001100101011111: color_data = 12'b111011101110;
20'b01001001100101100000: color_data = 12'b111011101110;
20'b01001001100101100001: color_data = 12'b111011101110;
20'b01001001100101100011: color_data = 12'b111011101110;
20'b01001001100101100100: color_data = 12'b111011101110;
20'b01001001100101100101: color_data = 12'b111011101110;
20'b01001001100101100110: color_data = 12'b111011101110;
20'b01001001100101100111: color_data = 12'b111011101110;
20'b01001001100101101110: color_data = 12'b111011101110;
20'b01001001100101101111: color_data = 12'b111011101110;
20'b01001001100101110000: color_data = 12'b111011101110;
20'b01001001100101110001: color_data = 12'b111011101110;
20'b01001001100101110010: color_data = 12'b111011101110;
20'b01001001100101110100: color_data = 12'b111111111111;
20'b01001001100101110101: color_data = 12'b111011101110;
20'b01001001100101110110: color_data = 12'b111011101110;
20'b01001001100101110111: color_data = 12'b111011101110;
20'b01001001100101111000: color_data = 12'b111011101110;
20'b01001001100110001010: color_data = 12'b111011101110;
20'b01001001100110001011: color_data = 12'b111011101110;
20'b01001001100110001100: color_data = 12'b111011101110;
20'b01001001100110001101: color_data = 12'b111011101110;
20'b01001001100110001110: color_data = 12'b111011101110;
20'b01001001100110010000: color_data = 12'b111011101110;
20'b01001001100110010001: color_data = 12'b111011101110;
20'b01001001100110010010: color_data = 12'b111011101110;
20'b01001001100110010011: color_data = 12'b111111111111;
20'b01001001110011110001: color_data = 12'b111011101110;
20'b01001001110011110010: color_data = 12'b111111111111;
20'b01001001110011110011: color_data = 12'b111011101110;
20'b01001001110011110100: color_data = 12'b111011101110;
20'b01001001110011110101: color_data = 12'b111011101110;
20'b01001001110011110111: color_data = 12'b111011101110;
20'b01001001110011111000: color_data = 12'b111011101110;
20'b01001001110011111001: color_data = 12'b111011101110;
20'b01001001110011111010: color_data = 12'b111011101110;
20'b01001001110011111100: color_data = 12'b111011101110;
20'b01001001110011111101: color_data = 12'b111011101110;
20'b01001001110011111110: color_data = 12'b111011101110;
20'b01001001110011111111: color_data = 12'b111011101110;
20'b01001001110100000000: color_data = 12'b111011101110;
20'b01001001110100000010: color_data = 12'b111011101110;
20'b01001001110100000011: color_data = 12'b111011101110;
20'b01001001110100000100: color_data = 12'b111011101110;
20'b01001001110100000101: color_data = 12'b111011101110;
20'b01001001110100000111: color_data = 12'b111011101110;
20'b01001001110100001000: color_data = 12'b111111111111;
20'b01001001110100001001: color_data = 12'b111011101110;
20'b01001001110100001010: color_data = 12'b111011101110;
20'b01001001110100001011: color_data = 12'b111111111111;
20'b01001001110100100010: color_data = 12'b111111111111;
20'b01001001110100100011: color_data = 12'b111011101110;
20'b01001001110100100100: color_data = 12'b111011101110;
20'b01001001110100100101: color_data = 12'b111011101110;
20'b01001001110100100110: color_data = 12'b111011101110;
20'b01001001110100101000: color_data = 12'b111011101110;
20'b01001001110100101001: color_data = 12'b111011101110;
20'b01001001110100101010: color_data = 12'b111011101110;
20'b01001001110100101011: color_data = 12'b111011101110;
20'b01001001110100101101: color_data = 12'b111011101110;
20'b01001001110100101110: color_data = 12'b111011101110;
20'b01001001110100101111: color_data = 12'b111011101110;
20'b01001001110100110000: color_data = 12'b111011101110;
20'b01001001110101000010: color_data = 12'b111011101110;
20'b01001001110101000011: color_data = 12'b111011101110;
20'b01001001110101000100: color_data = 12'b111011101110;
20'b01001001110101000101: color_data = 12'b111011101110;
20'b01001001110101000110: color_data = 12'b111011101110;
20'b01001001110101001000: color_data = 12'b111011101110;
20'b01001001110101001001: color_data = 12'b111011101110;
20'b01001001110101001010: color_data = 12'b111011101110;
20'b01001001110101001011: color_data = 12'b111111111111;
20'b01001001110101001100: color_data = 12'b111011101110;
20'b01001001110101001110: color_data = 12'b111111111111;
20'b01001001110101001111: color_data = 12'b111011101110;
20'b01001001110101010000: color_data = 12'b111011101110;
20'b01001001110101010001: color_data = 12'b111111111111;
20'b01001001110101010011: color_data = 12'b111011101110;
20'b01001001110101010100: color_data = 12'b111011101110;
20'b01001001110101010101: color_data = 12'b111011101110;
20'b01001001110101010110: color_data = 12'b111011101110;
20'b01001001110101011000: color_data = 12'b111011101110;
20'b01001001110101011001: color_data = 12'b111011101110;
20'b01001001110101011010: color_data = 12'b111011101110;
20'b01001001110101011011: color_data = 12'b111111111111;
20'b01001001110101011100: color_data = 12'b111011101110;
20'b01001001110101011110: color_data = 12'b111111111111;
20'b01001001110101011111: color_data = 12'b111011101110;
20'b01001001110101100000: color_data = 12'b111011101110;
20'b01001001110101100001: color_data = 12'b111111111111;
20'b01001001110101100011: color_data = 12'b111011101110;
20'b01001001110101100100: color_data = 12'b111111111111;
20'b01001001110101100101: color_data = 12'b111011101110;
20'b01001001110101100110: color_data = 12'b111011101110;
20'b01001001110101100111: color_data = 12'b111011101110;
20'b01001001110101101110: color_data = 12'b111111111111;
20'b01001001110101101111: color_data = 12'b111011101110;
20'b01001001110101110000: color_data = 12'b111011101110;
20'b01001001110101110001: color_data = 12'b111011101110;
20'b01001001110101110010: color_data = 12'b111011101110;
20'b01001001110101110100: color_data = 12'b111011101110;
20'b01001001110101110101: color_data = 12'b111011101110;
20'b01001001110101110110: color_data = 12'b111011101110;
20'b01001001110101110111: color_data = 12'b111011101110;
20'b01001001110101111000: color_data = 12'b111011101110;
20'b01001001110110001010: color_data = 12'b111111111111;
20'b01001001110110001011: color_data = 12'b111011101110;
20'b01001001110110001100: color_data = 12'b111011101110;
20'b01001001110110001101: color_data = 12'b111011101110;
20'b01001001110110001110: color_data = 12'b111011101110;
20'b01001001110110010000: color_data = 12'b111011101110;
20'b01001001110110010001: color_data = 12'b111011101110;
20'b01001001110110010010: color_data = 12'b111011101110;
20'b01001001110110010011: color_data = 12'b111011101110;
default: color_data = 12'b0;

	endcase
	end
endmodule