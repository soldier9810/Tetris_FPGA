`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/22/2025 04:19:03 PM
// Design Name: 
// Module Name: level1bmp_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// Dependencies: 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:

module level1bmp_rom
	(
		input clk,
		input [9:0] row,
		input [9:0] col,
		output reg [11:0] color_data,
		input ce
	);
	    (* rom_style = "block" *)
	
	reg [9:0] row_reg;
	reg [9:0] col_reg;
	always @(posedge clk)
		begin
		if (ce) begin
		row_reg <= row;
		col_reg <= col;
		end
		end
	always @(*) begin
	case ({row_reg, col_reg})
		20'b00010100010011010011: color_data = 12'b000000001111;
20'b00010100010011010100: color_data = 12'b000000001111;
20'b00010100010011010101: color_data = 12'b000000001111;
20'b00010100010011010110: color_data = 12'b000000001111;
20'b00010100010011010111: color_data = 12'b000000001111;
20'b00010100010011011000: color_data = 12'b000000001111;
20'b00010100010011011001: color_data = 12'b000000001111;
20'b00010100010011011010: color_data = 12'b000000001111;
20'b00010100010011011011: color_data = 12'b000000001111;
20'b00010100010011011100: color_data = 12'b000000001111;
20'b00010100010011011101: color_data = 12'b000000001111;
20'b00010100010011011110: color_data = 12'b000000001111;
20'b00010100010011011111: color_data = 12'b000000001111;
20'b00010100010011100000: color_data = 12'b000000001111;
20'b00010100010011100001: color_data = 12'b000000001111;
20'b00010100010011100010: color_data = 12'b000000001111;
20'b00010100010011100011: color_data = 12'b000000001111;
20'b00010100010011100100: color_data = 12'b000000001111;
20'b00010100010011100101: color_data = 12'b000000001111;
20'b00010100010011100110: color_data = 12'b000000001111;
20'b00010100010011100111: color_data = 12'b000000001111;
20'b00010100010011101000: color_data = 12'b000000001111;
20'b00010100010011101001: color_data = 12'b000000001111;
20'b00010100010011101010: color_data = 12'b000000001111;
20'b00010100010011101011: color_data = 12'b000000001111;
20'b00010100010011101100: color_data = 12'b000000001111;
20'b00010100010011101101: color_data = 12'b000000001111;
20'b00010100010011101110: color_data = 12'b000000001111;
20'b00010100010011101111: color_data = 12'b000000001111;
20'b00010100010011110000: color_data = 12'b000000001111;
20'b00010100010011110001: color_data = 12'b000000001111;
20'b00010100010011110010: color_data = 12'b000000001111;
20'b00010100010011110011: color_data = 12'b000000001111;
20'b00010100010011110100: color_data = 12'b000000001111;
20'b00010100010011110101: color_data = 12'b000000001111;
20'b00010100010011110110: color_data = 12'b000000001111;
20'b00010100010011110111: color_data = 12'b000000001111;
20'b00010100010011111000: color_data = 12'b000000001111;
20'b00010100010011111001: color_data = 12'b000000001111;
20'b00010100010011111010: color_data = 12'b000000001111;
20'b00010100010011111011: color_data = 12'b000000001111;
20'b00010100010100000101: color_data = 12'b000001101111;
20'b00010100010100000110: color_data = 12'b000001101111;
20'b00010100010100000111: color_data = 12'b000001101111;
20'b00010100010100001000: color_data = 12'b000001101111;
20'b00010100010100001001: color_data = 12'b000001101111;
20'b00010100010100001010: color_data = 12'b000001101111;
20'b00010100010100001011: color_data = 12'b000001101111;
20'b00010100010100001100: color_data = 12'b000001101111;
20'b00010100010100001101: color_data = 12'b000001101111;
20'b00010100010100001110: color_data = 12'b000001101111;
20'b00010100010100001111: color_data = 12'b000001101111;
20'b00010100010100010000: color_data = 12'b000001101111;
20'b00010100010100010001: color_data = 12'b000001101111;
20'b00010100010100010010: color_data = 12'b000001101111;
20'b00010100010100010011: color_data = 12'b000001101111;
20'b00010100010100010100: color_data = 12'b000001101111;
20'b00010100010100010101: color_data = 12'b000001101111;
20'b00010100010100010110: color_data = 12'b000001101111;
20'b00010100010100010111: color_data = 12'b000001101111;
20'b00010100010100011000: color_data = 12'b000001101111;
20'b00010100010100011001: color_data = 12'b000001101111;
20'b00010100010100011010: color_data = 12'b000001101111;
20'b00010100010100011011: color_data = 12'b000001101111;
20'b00010100010100011100: color_data = 12'b000001101111;
20'b00010100010100011101: color_data = 12'b000001101111;
20'b00010100010100011110: color_data = 12'b000001101111;
20'b00010100010100011111: color_data = 12'b000001101111;
20'b00010100010100100000: color_data = 12'b000001101111;
20'b00010100010100100001: color_data = 12'b000001101111;
20'b00010100010100100010: color_data = 12'b000001101111;
20'b00010100010100100011: color_data = 12'b000001101111;
20'b00010100010100100100: color_data = 12'b000001101111;
20'b00010100010100101101: color_data = 12'b000011111111;
20'b00010100010100101110: color_data = 12'b000011111111;
20'b00010100010100101111: color_data = 12'b000011111111;
20'b00010100010100110000: color_data = 12'b000011111111;
20'b00010100010100110001: color_data = 12'b000011111111;
20'b00010100010100110010: color_data = 12'b000011111111;
20'b00010100010100110011: color_data = 12'b000011111111;
20'b00010100010100110100: color_data = 12'b000011111111;
20'b00010100010100110101: color_data = 12'b000011111111;
20'b00010100010100110110: color_data = 12'b000011111111;
20'b00010100010100110111: color_data = 12'b000011111111;
20'b00010100010100111000: color_data = 12'b000011111111;
20'b00010100010100111001: color_data = 12'b000011111111;
20'b00010100010100111010: color_data = 12'b000011111111;
20'b00010100010100111011: color_data = 12'b000011111111;
20'b00010100010100111100: color_data = 12'b000011111111;
20'b00010100010100111101: color_data = 12'b000011111111;
20'b00010100010100111110: color_data = 12'b000011111111;
20'b00010100010100111111: color_data = 12'b000011111111;
20'b00010100010101000000: color_data = 12'b000011111111;
20'b00010100010101000001: color_data = 12'b000011111111;
20'b00010100010101000010: color_data = 12'b000011111111;
20'b00010100010101000011: color_data = 12'b000011111111;
20'b00010100010101000100: color_data = 12'b000011111111;
20'b00010100010101000101: color_data = 12'b000011111111;
20'b00010100010101000110: color_data = 12'b000011111111;
20'b00010100010101000111: color_data = 12'b000011111111;
20'b00010100010101001000: color_data = 12'b000011111111;
20'b00010100010101001001: color_data = 12'b000011111111;
20'b00010100010101001010: color_data = 12'b000011111111;
20'b00010100010101001011: color_data = 12'b000011111111;
20'b00010100010101001100: color_data = 12'b000011111111;
20'b00010100010101001101: color_data = 12'b000011111111;
20'b00010100010101001110: color_data = 12'b000011111111;
20'b00010100010101001111: color_data = 12'b000011111111;
20'b00010100010101010000: color_data = 12'b000011111111;
20'b00010100010101010001: color_data = 12'b000011111111;
20'b00010100010101010010: color_data = 12'b000011111111;
20'b00010100010101010011: color_data = 12'b000011111111;
20'b00010100010101010100: color_data = 12'b000011111111;
20'b00010100010101010101: color_data = 12'b000011111111;
20'b00010100010101011111: color_data = 12'b111101110000;
20'b00010100010101100000: color_data = 12'b111101110000;
20'b00010100010101100001: color_data = 12'b111101110000;
20'b00010100010101100010: color_data = 12'b111101110000;
20'b00010100010101100011: color_data = 12'b111101110000;
20'b00010100010101100100: color_data = 12'b111101110000;
20'b00010100010101100101: color_data = 12'b111101110000;
20'b00010100010101100110: color_data = 12'b111101110000;
20'b00010100010101100111: color_data = 12'b111101110000;
20'b00010100010101101000: color_data = 12'b111101110000;
20'b00010100010101101001: color_data = 12'b111101110000;
20'b00010100010101101010: color_data = 12'b111101110000;
20'b00010100010101101011: color_data = 12'b111101110000;
20'b00010100010101101100: color_data = 12'b111101110000;
20'b00010100010101101101: color_data = 12'b111101110000;
20'b00010100010101101110: color_data = 12'b111101110000;
20'b00010100010101101111: color_data = 12'b111101110000;
20'b00010100010101110000: color_data = 12'b111101110000;
20'b00010100010101110001: color_data = 12'b111101110000;
20'b00010100010101110010: color_data = 12'b111101110000;
20'b00010100010101110011: color_data = 12'b111101110000;
20'b00010100010101110100: color_data = 12'b111101110000;
20'b00010100010101110101: color_data = 12'b111101110000;
20'b00010100010101110110: color_data = 12'b111101110000;
20'b00010100010101110111: color_data = 12'b111101110000;
20'b00010100010101111000: color_data = 12'b111101110000;
20'b00010100010101111001: color_data = 12'b111101110000;
20'b00010100010101111010: color_data = 12'b111101110000;
20'b00010100010101111011: color_data = 12'b111101110000;
20'b00010100010101111100: color_data = 12'b111101110000;
20'b00010100010101111101: color_data = 12'b111101110000;
20'b00010100010101111110: color_data = 12'b111101110000;
20'b00010100010110000111: color_data = 12'b000011110000;
20'b00010100010110001000: color_data = 12'b000011110000;
20'b00010100010110001001: color_data = 12'b000011110000;
20'b00010100010110001010: color_data = 12'b000011110000;
20'b00010100010110001011: color_data = 12'b000011110000;
20'b00010100010110001100: color_data = 12'b000011110000;
20'b00010100010110001101: color_data = 12'b000011110000;
20'b00010100010110001110: color_data = 12'b000011110000;
20'b00010100010110001111: color_data = 12'b000011110000;
20'b00010100010110011000: color_data = 12'b111100001111;
20'b00010100010110011001: color_data = 12'b111100001111;
20'b00010100010110011010: color_data = 12'b111100001111;
20'b00010100010110011011: color_data = 12'b111100001111;
20'b00010100010110011100: color_data = 12'b111100001111;
20'b00010100010110011101: color_data = 12'b111100001111;
20'b00010100010110011110: color_data = 12'b111100001111;
20'b00010100010110011111: color_data = 12'b111100001111;
20'b00010100010110100000: color_data = 12'b111100001111;
20'b00010100010110100001: color_data = 12'b111100001111;
20'b00010100010110100010: color_data = 12'b111100001111;
20'b00010100010110100011: color_data = 12'b111100001111;
20'b00010100010110100100: color_data = 12'b111100001111;
20'b00010100010110100101: color_data = 12'b111100001111;
20'b00010100010110100110: color_data = 12'b111100001111;
20'b00010100010110100111: color_data = 12'b111100001111;
20'b00010100010110101000: color_data = 12'b111100001111;
20'b00010100010110101001: color_data = 12'b111100001111;
20'b00010100010110101010: color_data = 12'b111100001111;
20'b00010100010110101011: color_data = 12'b111100001111;
20'b00010100010110101100: color_data = 12'b111100001111;
20'b00010100010110101101: color_data = 12'b111100001111;
20'b00010100010110101110: color_data = 12'b111100001111;
20'b00010100010110101111: color_data = 12'b111100001111;
20'b00010100010110110000: color_data = 12'b111100001111;
20'b00010100010110110001: color_data = 12'b111100001111;
20'b00010100010110110010: color_data = 12'b111100001111;
20'b00010100010110110011: color_data = 12'b111100001111;
20'b00010100010110110100: color_data = 12'b111100001111;
20'b00010100010110110101: color_data = 12'b111100001111;
20'b00010100010110110110: color_data = 12'b111100001111;
20'b00010100010110110111: color_data = 12'b111100001111;
20'b00010100100011010011: color_data = 12'b000000001111;
20'b00010100100011010100: color_data = 12'b000000001111;
20'b00010100100011010101: color_data = 12'b000000001111;
20'b00010100100011010110: color_data = 12'b000000001111;
20'b00010100100011010111: color_data = 12'b000000001111;
20'b00010100100011011000: color_data = 12'b000000001111;
20'b00010100100011011001: color_data = 12'b000000001111;
20'b00010100100011011010: color_data = 12'b000000001111;
20'b00010100100011011011: color_data = 12'b000000001111;
20'b00010100100011011100: color_data = 12'b000000001111;
20'b00010100100011011101: color_data = 12'b000000001111;
20'b00010100100011011110: color_data = 12'b000000001111;
20'b00010100100011011111: color_data = 12'b000000001111;
20'b00010100100011100000: color_data = 12'b000000001111;
20'b00010100100011100001: color_data = 12'b000000001111;
20'b00010100100011100010: color_data = 12'b000000001111;
20'b00010100100011100011: color_data = 12'b000000001111;
20'b00010100100011100100: color_data = 12'b000000001111;
20'b00010100100011100101: color_data = 12'b000000001111;
20'b00010100100011100110: color_data = 12'b000000001111;
20'b00010100100011100111: color_data = 12'b000000001111;
20'b00010100100011101000: color_data = 12'b000000001111;
20'b00010100100011101001: color_data = 12'b000000001111;
20'b00010100100011101010: color_data = 12'b000000001111;
20'b00010100100011101011: color_data = 12'b000000001111;
20'b00010100100011101100: color_data = 12'b000000001111;
20'b00010100100011101101: color_data = 12'b000000001111;
20'b00010100100011101110: color_data = 12'b000000001111;
20'b00010100100011101111: color_data = 12'b000000001111;
20'b00010100100011110000: color_data = 12'b000000001111;
20'b00010100100011110001: color_data = 12'b000000001111;
20'b00010100100011110010: color_data = 12'b000000001111;
20'b00010100100011110011: color_data = 12'b000000001111;
20'b00010100100011110100: color_data = 12'b000000001111;
20'b00010100100011110101: color_data = 12'b000000001111;
20'b00010100100011110110: color_data = 12'b000000001111;
20'b00010100100011110111: color_data = 12'b000000001111;
20'b00010100100011111000: color_data = 12'b000000001111;
20'b00010100100011111001: color_data = 12'b000000001111;
20'b00010100100011111010: color_data = 12'b000000001111;
20'b00010100100011111011: color_data = 12'b000000001111;
20'b00010100100100000101: color_data = 12'b000001101111;
20'b00010100100100000110: color_data = 12'b000001101111;
20'b00010100100100000111: color_data = 12'b000001101111;
20'b00010100100100001000: color_data = 12'b000001101111;
20'b00010100100100001001: color_data = 12'b000001101111;
20'b00010100100100001010: color_data = 12'b000001101111;
20'b00010100100100001011: color_data = 12'b000001101111;
20'b00010100100100001100: color_data = 12'b000001101111;
20'b00010100100100001101: color_data = 12'b000001101111;
20'b00010100100100001110: color_data = 12'b000001101111;
20'b00010100100100001111: color_data = 12'b000001101111;
20'b00010100100100010000: color_data = 12'b000001101111;
20'b00010100100100010001: color_data = 12'b000001101111;
20'b00010100100100010010: color_data = 12'b000001101111;
20'b00010100100100010011: color_data = 12'b000001101111;
20'b00010100100100010100: color_data = 12'b000001101111;
20'b00010100100100010101: color_data = 12'b000001101111;
20'b00010100100100010110: color_data = 12'b000001101111;
20'b00010100100100010111: color_data = 12'b000001101111;
20'b00010100100100011000: color_data = 12'b000001101111;
20'b00010100100100011001: color_data = 12'b000001101111;
20'b00010100100100011010: color_data = 12'b000001101111;
20'b00010100100100011011: color_data = 12'b000001101111;
20'b00010100100100011100: color_data = 12'b000001101111;
20'b00010100100100011101: color_data = 12'b000001101111;
20'b00010100100100011110: color_data = 12'b000001101111;
20'b00010100100100011111: color_data = 12'b000001101111;
20'b00010100100100100000: color_data = 12'b000001101111;
20'b00010100100100100001: color_data = 12'b000001101111;
20'b00010100100100100010: color_data = 12'b000001101111;
20'b00010100100100100011: color_data = 12'b000001101111;
20'b00010100100100100100: color_data = 12'b000001101111;
20'b00010100100100101101: color_data = 12'b000011111111;
20'b00010100100100101110: color_data = 12'b000011111111;
20'b00010100100100101111: color_data = 12'b000011111111;
20'b00010100100100110000: color_data = 12'b000011111111;
20'b00010100100100110001: color_data = 12'b000011111111;
20'b00010100100100110010: color_data = 12'b000011111111;
20'b00010100100100110011: color_data = 12'b000011111111;
20'b00010100100100110100: color_data = 12'b000011111111;
20'b00010100100100110101: color_data = 12'b000011111111;
20'b00010100100100110110: color_data = 12'b000011111111;
20'b00010100100100110111: color_data = 12'b000011111111;
20'b00010100100100111000: color_data = 12'b000011111111;
20'b00010100100100111001: color_data = 12'b000011111111;
20'b00010100100100111010: color_data = 12'b000011111111;
20'b00010100100100111011: color_data = 12'b000011111111;
20'b00010100100100111100: color_data = 12'b000011111111;
20'b00010100100100111101: color_data = 12'b000011111111;
20'b00010100100100111110: color_data = 12'b000011111111;
20'b00010100100100111111: color_data = 12'b000011111111;
20'b00010100100101000000: color_data = 12'b000011111111;
20'b00010100100101000001: color_data = 12'b000011111111;
20'b00010100100101000010: color_data = 12'b000011111111;
20'b00010100100101000011: color_data = 12'b000011111111;
20'b00010100100101000100: color_data = 12'b000011111111;
20'b00010100100101000101: color_data = 12'b000011111111;
20'b00010100100101000110: color_data = 12'b000011111111;
20'b00010100100101000111: color_data = 12'b000011111111;
20'b00010100100101001000: color_data = 12'b000011111111;
20'b00010100100101001001: color_data = 12'b000011111111;
20'b00010100100101001010: color_data = 12'b000011111111;
20'b00010100100101001011: color_data = 12'b000011111111;
20'b00010100100101001100: color_data = 12'b000011111111;
20'b00010100100101001101: color_data = 12'b000011111111;
20'b00010100100101001110: color_data = 12'b000011111111;
20'b00010100100101001111: color_data = 12'b000011111111;
20'b00010100100101010000: color_data = 12'b000011111111;
20'b00010100100101010001: color_data = 12'b000011111111;
20'b00010100100101010010: color_data = 12'b000011111111;
20'b00010100100101010011: color_data = 12'b000011111111;
20'b00010100100101010100: color_data = 12'b000011111111;
20'b00010100100101010101: color_data = 12'b000011111111;
20'b00010100100101011111: color_data = 12'b111101110000;
20'b00010100100101100000: color_data = 12'b111101110000;
20'b00010100100101100001: color_data = 12'b111101110000;
20'b00010100100101100010: color_data = 12'b111101110000;
20'b00010100100101100011: color_data = 12'b111101110000;
20'b00010100100101100100: color_data = 12'b111101110000;
20'b00010100100101100101: color_data = 12'b111101110000;
20'b00010100100101100110: color_data = 12'b111101110000;
20'b00010100100101100111: color_data = 12'b111101110000;
20'b00010100100101101000: color_data = 12'b111101110000;
20'b00010100100101101001: color_data = 12'b111101110000;
20'b00010100100101101010: color_data = 12'b111101110000;
20'b00010100100101101011: color_data = 12'b111101110000;
20'b00010100100101101100: color_data = 12'b111101110000;
20'b00010100100101101101: color_data = 12'b111101110000;
20'b00010100100101101110: color_data = 12'b111101110000;
20'b00010100100101101111: color_data = 12'b111101110000;
20'b00010100100101110000: color_data = 12'b111101110000;
20'b00010100100101110001: color_data = 12'b111101110000;
20'b00010100100101110010: color_data = 12'b111101110000;
20'b00010100100101110011: color_data = 12'b111101110000;
20'b00010100100101110100: color_data = 12'b111101110000;
20'b00010100100101110101: color_data = 12'b111101110000;
20'b00010100100101110110: color_data = 12'b111101110000;
20'b00010100100101110111: color_data = 12'b111101110000;
20'b00010100100101111000: color_data = 12'b111101110000;
20'b00010100100101111001: color_data = 12'b111101110000;
20'b00010100100101111010: color_data = 12'b111101110000;
20'b00010100100101111011: color_data = 12'b111101110000;
20'b00010100100101111100: color_data = 12'b111101110000;
20'b00010100100101111101: color_data = 12'b111101110000;
20'b00010100100101111110: color_data = 12'b111101110000;
20'b00010100100110000111: color_data = 12'b000011110000;
20'b00010100100110001000: color_data = 12'b000011110000;
20'b00010100100110001001: color_data = 12'b000011110000;
20'b00010100100110001010: color_data = 12'b000011110000;
20'b00010100100110001011: color_data = 12'b000011110000;
20'b00010100100110001100: color_data = 12'b000011110000;
20'b00010100100110001101: color_data = 12'b000011110000;
20'b00010100100110001110: color_data = 12'b000011110000;
20'b00010100100110001111: color_data = 12'b000011110000;
20'b00010100100110011000: color_data = 12'b111100001111;
20'b00010100100110011001: color_data = 12'b111100001111;
20'b00010100100110011010: color_data = 12'b111100001111;
20'b00010100100110011011: color_data = 12'b111100001111;
20'b00010100100110011100: color_data = 12'b111100001111;
20'b00010100100110011101: color_data = 12'b111100001111;
20'b00010100100110011110: color_data = 12'b111100001111;
20'b00010100100110011111: color_data = 12'b111100001111;
20'b00010100100110100000: color_data = 12'b111100001111;
20'b00010100100110100001: color_data = 12'b111100001111;
20'b00010100100110100010: color_data = 12'b111100001111;
20'b00010100100110100011: color_data = 12'b111100001111;
20'b00010100100110100100: color_data = 12'b111100001111;
20'b00010100100110100101: color_data = 12'b111100001111;
20'b00010100100110100110: color_data = 12'b111100001111;
20'b00010100100110100111: color_data = 12'b111100001111;
20'b00010100100110101000: color_data = 12'b111100001111;
20'b00010100100110101001: color_data = 12'b111100001111;
20'b00010100100110101010: color_data = 12'b111100001111;
20'b00010100100110101011: color_data = 12'b111100001111;
20'b00010100100110101100: color_data = 12'b111100001111;
20'b00010100100110101101: color_data = 12'b111100001111;
20'b00010100100110101110: color_data = 12'b111100001111;
20'b00010100100110101111: color_data = 12'b111100001111;
20'b00010100100110110000: color_data = 12'b111100001111;
20'b00010100100110110001: color_data = 12'b111100001111;
20'b00010100100110110010: color_data = 12'b111100001111;
20'b00010100100110110011: color_data = 12'b111100001111;
20'b00010100100110110100: color_data = 12'b111100001111;
20'b00010100100110110101: color_data = 12'b111100001111;
20'b00010100100110110110: color_data = 12'b111100001111;
20'b00010100100110110111: color_data = 12'b111100001111;
20'b00010100110011010011: color_data = 12'b000000001111;
20'b00010100110011010100: color_data = 12'b000000001111;
20'b00010100110011010101: color_data = 12'b000000001111;
20'b00010100110011010110: color_data = 12'b000000001111;
20'b00010100110011010111: color_data = 12'b000000001111;
20'b00010100110011011000: color_data = 12'b000000001111;
20'b00010100110011011001: color_data = 12'b000000001111;
20'b00010100110011011010: color_data = 12'b000000001111;
20'b00010100110011011011: color_data = 12'b000000001111;
20'b00010100110011011100: color_data = 12'b000000001111;
20'b00010100110011011101: color_data = 12'b000000001111;
20'b00010100110011011110: color_data = 12'b000000001111;
20'b00010100110011011111: color_data = 12'b000000001111;
20'b00010100110011100000: color_data = 12'b000000001111;
20'b00010100110011100001: color_data = 12'b000000001111;
20'b00010100110011100010: color_data = 12'b000000001111;
20'b00010100110011100011: color_data = 12'b000000001111;
20'b00010100110011100100: color_data = 12'b000000001111;
20'b00010100110011100101: color_data = 12'b000000001111;
20'b00010100110011100110: color_data = 12'b000000001111;
20'b00010100110011100111: color_data = 12'b000000001111;
20'b00010100110011101000: color_data = 12'b000000001111;
20'b00010100110011101001: color_data = 12'b000000001111;
20'b00010100110011101010: color_data = 12'b000000001111;
20'b00010100110011101011: color_data = 12'b000000001111;
20'b00010100110011101100: color_data = 12'b000000001111;
20'b00010100110011101101: color_data = 12'b000000001111;
20'b00010100110011101110: color_data = 12'b000000001111;
20'b00010100110011101111: color_data = 12'b000000001111;
20'b00010100110011110000: color_data = 12'b000000001111;
20'b00010100110011110001: color_data = 12'b000000001111;
20'b00010100110011110010: color_data = 12'b000000001111;
20'b00010100110011110011: color_data = 12'b000000001111;
20'b00010100110011110100: color_data = 12'b000000001111;
20'b00010100110011110101: color_data = 12'b000000001111;
20'b00010100110011110110: color_data = 12'b000000001111;
20'b00010100110011110111: color_data = 12'b000000001111;
20'b00010100110011111000: color_data = 12'b000000001111;
20'b00010100110011111001: color_data = 12'b000000001111;
20'b00010100110011111010: color_data = 12'b000000001111;
20'b00010100110011111011: color_data = 12'b000000001111;
20'b00010100110100000101: color_data = 12'b000001101111;
20'b00010100110100000110: color_data = 12'b000001101111;
20'b00010100110100000111: color_data = 12'b000001101111;
20'b00010100110100001000: color_data = 12'b000001101111;
20'b00010100110100001001: color_data = 12'b000001101111;
20'b00010100110100001010: color_data = 12'b000001101111;
20'b00010100110100001011: color_data = 12'b000001101111;
20'b00010100110100001100: color_data = 12'b000001101111;
20'b00010100110100001101: color_data = 12'b000001101111;
20'b00010100110100001110: color_data = 12'b000001101111;
20'b00010100110100001111: color_data = 12'b000001101111;
20'b00010100110100010000: color_data = 12'b000001101111;
20'b00010100110100010001: color_data = 12'b000001101111;
20'b00010100110100010010: color_data = 12'b000001101111;
20'b00010100110100010011: color_data = 12'b000001101111;
20'b00010100110100010100: color_data = 12'b000001101111;
20'b00010100110100010101: color_data = 12'b000001101111;
20'b00010100110100010110: color_data = 12'b000001101111;
20'b00010100110100010111: color_data = 12'b000001101111;
20'b00010100110100011000: color_data = 12'b000001101111;
20'b00010100110100011001: color_data = 12'b000001101111;
20'b00010100110100011010: color_data = 12'b000001101111;
20'b00010100110100011011: color_data = 12'b000001101111;
20'b00010100110100011100: color_data = 12'b000001101111;
20'b00010100110100011101: color_data = 12'b000001101111;
20'b00010100110100011110: color_data = 12'b000001101111;
20'b00010100110100011111: color_data = 12'b000001101111;
20'b00010100110100100000: color_data = 12'b000001101111;
20'b00010100110100100001: color_data = 12'b000001101111;
20'b00010100110100100010: color_data = 12'b000001101111;
20'b00010100110100100011: color_data = 12'b000001101111;
20'b00010100110100100100: color_data = 12'b000001101111;
20'b00010100110100101101: color_data = 12'b000011111111;
20'b00010100110100101110: color_data = 12'b000011111111;
20'b00010100110100101111: color_data = 12'b000011111111;
20'b00010100110100110000: color_data = 12'b000011111111;
20'b00010100110100110001: color_data = 12'b000011111111;
20'b00010100110100110010: color_data = 12'b000011111111;
20'b00010100110100110011: color_data = 12'b000011111111;
20'b00010100110100110100: color_data = 12'b000011111111;
20'b00010100110100110101: color_data = 12'b000011111111;
20'b00010100110100110110: color_data = 12'b000011111111;
20'b00010100110100110111: color_data = 12'b000011111111;
20'b00010100110100111000: color_data = 12'b000011111111;
20'b00010100110100111001: color_data = 12'b000011111111;
20'b00010100110100111010: color_data = 12'b000011111111;
20'b00010100110100111011: color_data = 12'b000011111111;
20'b00010100110100111100: color_data = 12'b000011111111;
20'b00010100110100111101: color_data = 12'b000011111111;
20'b00010100110100111110: color_data = 12'b000011111111;
20'b00010100110100111111: color_data = 12'b000011111111;
20'b00010100110101000000: color_data = 12'b000011111111;
20'b00010100110101000001: color_data = 12'b000011111111;
20'b00010100110101000010: color_data = 12'b000011111111;
20'b00010100110101000011: color_data = 12'b000011111111;
20'b00010100110101000100: color_data = 12'b000011111111;
20'b00010100110101000101: color_data = 12'b000011111111;
20'b00010100110101000110: color_data = 12'b000011111111;
20'b00010100110101000111: color_data = 12'b000011111111;
20'b00010100110101001000: color_data = 12'b000011111111;
20'b00010100110101001001: color_data = 12'b000011111111;
20'b00010100110101001010: color_data = 12'b000011111111;
20'b00010100110101001011: color_data = 12'b000011111111;
20'b00010100110101001100: color_data = 12'b000011111111;
20'b00010100110101001101: color_data = 12'b000011111111;
20'b00010100110101001110: color_data = 12'b000011111111;
20'b00010100110101001111: color_data = 12'b000011111111;
20'b00010100110101010000: color_data = 12'b000011111111;
20'b00010100110101010001: color_data = 12'b000011111111;
20'b00010100110101010010: color_data = 12'b000011111111;
20'b00010100110101010011: color_data = 12'b000011111111;
20'b00010100110101010100: color_data = 12'b000011111111;
20'b00010100110101010101: color_data = 12'b000011111111;
20'b00010100110101011111: color_data = 12'b111101110000;
20'b00010100110101100000: color_data = 12'b111101110000;
20'b00010100110101100001: color_data = 12'b111101110000;
20'b00010100110101100010: color_data = 12'b111101110000;
20'b00010100110101100011: color_data = 12'b111101110000;
20'b00010100110101100100: color_data = 12'b111101110000;
20'b00010100110101100101: color_data = 12'b111101110000;
20'b00010100110101100110: color_data = 12'b111101110000;
20'b00010100110101100111: color_data = 12'b111101110000;
20'b00010100110101101000: color_data = 12'b111101110000;
20'b00010100110101101001: color_data = 12'b111101110000;
20'b00010100110101101010: color_data = 12'b111101110000;
20'b00010100110101101011: color_data = 12'b111101110000;
20'b00010100110101101100: color_data = 12'b111101110000;
20'b00010100110101101101: color_data = 12'b111101110000;
20'b00010100110101101110: color_data = 12'b111101110000;
20'b00010100110101101111: color_data = 12'b111101110000;
20'b00010100110101110000: color_data = 12'b111101110000;
20'b00010100110101110001: color_data = 12'b111101110000;
20'b00010100110101110010: color_data = 12'b111101110000;
20'b00010100110101110011: color_data = 12'b111101110000;
20'b00010100110101110100: color_data = 12'b111101110000;
20'b00010100110101110101: color_data = 12'b111101110000;
20'b00010100110101110110: color_data = 12'b111101110000;
20'b00010100110101110111: color_data = 12'b111101110000;
20'b00010100110101111000: color_data = 12'b111101110000;
20'b00010100110101111001: color_data = 12'b111101110000;
20'b00010100110101111010: color_data = 12'b111101110000;
20'b00010100110101111011: color_data = 12'b111101110000;
20'b00010100110101111100: color_data = 12'b111101110000;
20'b00010100110101111101: color_data = 12'b111101110000;
20'b00010100110101111110: color_data = 12'b111101110000;
20'b00010100110110000111: color_data = 12'b000011110000;
20'b00010100110110001000: color_data = 12'b000011110000;
20'b00010100110110001001: color_data = 12'b000011110000;
20'b00010100110110001010: color_data = 12'b000011110000;
20'b00010100110110001011: color_data = 12'b000011110000;
20'b00010100110110001100: color_data = 12'b000011110000;
20'b00010100110110001101: color_data = 12'b000011110000;
20'b00010100110110001110: color_data = 12'b000011110000;
20'b00010100110110001111: color_data = 12'b000011110000;
20'b00010100110110011000: color_data = 12'b111100001111;
20'b00010100110110011001: color_data = 12'b111100001111;
20'b00010100110110011010: color_data = 12'b111100001111;
20'b00010100110110011011: color_data = 12'b111100001111;
20'b00010100110110011100: color_data = 12'b111100001111;
20'b00010100110110011101: color_data = 12'b111100001111;
20'b00010100110110011110: color_data = 12'b111100001111;
20'b00010100110110011111: color_data = 12'b111100001111;
20'b00010100110110100000: color_data = 12'b111100001111;
20'b00010100110110100001: color_data = 12'b111100001111;
20'b00010100110110100010: color_data = 12'b111100001111;
20'b00010100110110100011: color_data = 12'b111100001111;
20'b00010100110110100100: color_data = 12'b111100001111;
20'b00010100110110100101: color_data = 12'b111100001111;
20'b00010100110110100110: color_data = 12'b111100001111;
20'b00010100110110100111: color_data = 12'b111100001111;
20'b00010100110110101000: color_data = 12'b111100001111;
20'b00010100110110101001: color_data = 12'b111100001111;
20'b00010100110110101010: color_data = 12'b111100001111;
20'b00010100110110101011: color_data = 12'b111100001111;
20'b00010100110110101100: color_data = 12'b111100001111;
20'b00010100110110101101: color_data = 12'b111100001111;
20'b00010100110110101110: color_data = 12'b111100001111;
20'b00010100110110101111: color_data = 12'b111100001111;
20'b00010100110110110000: color_data = 12'b111100001111;
20'b00010100110110110001: color_data = 12'b111100001111;
20'b00010100110110110010: color_data = 12'b111100001111;
20'b00010100110110110011: color_data = 12'b111100001111;
20'b00010100110110110100: color_data = 12'b111100001111;
20'b00010100110110110101: color_data = 12'b111100001111;
20'b00010100110110110110: color_data = 12'b111100001111;
20'b00010100110110110111: color_data = 12'b111100001111;
20'b00010101000011010011: color_data = 12'b000000001111;
20'b00010101000011010100: color_data = 12'b000000001111;
20'b00010101000011010101: color_data = 12'b000000001111;
20'b00010101000011010110: color_data = 12'b000000001111;
20'b00010101000011010111: color_data = 12'b000000001111;
20'b00010101000011011000: color_data = 12'b000000001111;
20'b00010101000011011001: color_data = 12'b000000001111;
20'b00010101000011011010: color_data = 12'b000000001111;
20'b00010101000011011011: color_data = 12'b000000001111;
20'b00010101000011011100: color_data = 12'b000000001111;
20'b00010101000011011101: color_data = 12'b000000001111;
20'b00010101000011011110: color_data = 12'b000000001111;
20'b00010101000011011111: color_data = 12'b000000001111;
20'b00010101000011100000: color_data = 12'b000000001111;
20'b00010101000011100001: color_data = 12'b000000001111;
20'b00010101000011100010: color_data = 12'b000000001111;
20'b00010101000011100011: color_data = 12'b000000001111;
20'b00010101000011100100: color_data = 12'b000000001111;
20'b00010101000011100101: color_data = 12'b000000001111;
20'b00010101000011100110: color_data = 12'b000000001111;
20'b00010101000011100111: color_data = 12'b000000001111;
20'b00010101000011101000: color_data = 12'b000000001111;
20'b00010101000011101001: color_data = 12'b000000001111;
20'b00010101000011101010: color_data = 12'b000000001111;
20'b00010101000011101011: color_data = 12'b000000001111;
20'b00010101000011101100: color_data = 12'b000000001111;
20'b00010101000011101101: color_data = 12'b000000001111;
20'b00010101000011101110: color_data = 12'b000000001111;
20'b00010101000011101111: color_data = 12'b000000001111;
20'b00010101000011110000: color_data = 12'b000000001111;
20'b00010101000011110001: color_data = 12'b000000001111;
20'b00010101000011110010: color_data = 12'b000000001111;
20'b00010101000011110011: color_data = 12'b000000001111;
20'b00010101000011110100: color_data = 12'b000000001111;
20'b00010101000011110101: color_data = 12'b000000001111;
20'b00010101000011110110: color_data = 12'b000000001111;
20'b00010101000011110111: color_data = 12'b000000001111;
20'b00010101000011111000: color_data = 12'b000000001111;
20'b00010101000011111001: color_data = 12'b000000001111;
20'b00010101000011111010: color_data = 12'b000000001111;
20'b00010101000011111011: color_data = 12'b000000001111;
20'b00010101000100000101: color_data = 12'b000001101111;
20'b00010101000100000110: color_data = 12'b000001101111;
20'b00010101000100000111: color_data = 12'b000001101111;
20'b00010101000100001000: color_data = 12'b000001101111;
20'b00010101000100001001: color_data = 12'b000001101111;
20'b00010101000100001010: color_data = 12'b000001101111;
20'b00010101000100001011: color_data = 12'b000001101111;
20'b00010101000100001100: color_data = 12'b000001101111;
20'b00010101000100001101: color_data = 12'b000001101111;
20'b00010101000100001110: color_data = 12'b000001101111;
20'b00010101000100001111: color_data = 12'b000001101111;
20'b00010101000100010000: color_data = 12'b000001101111;
20'b00010101000100010001: color_data = 12'b000001101111;
20'b00010101000100010010: color_data = 12'b000001101111;
20'b00010101000100010011: color_data = 12'b000001101111;
20'b00010101000100010100: color_data = 12'b000001101111;
20'b00010101000100010101: color_data = 12'b000001101111;
20'b00010101000100010110: color_data = 12'b000001101111;
20'b00010101000100010111: color_data = 12'b000001101111;
20'b00010101000100011000: color_data = 12'b000001101111;
20'b00010101000100011001: color_data = 12'b000001101111;
20'b00010101000100011010: color_data = 12'b000001101111;
20'b00010101000100011011: color_data = 12'b000001101111;
20'b00010101000100011100: color_data = 12'b000001101111;
20'b00010101000100011101: color_data = 12'b000001101111;
20'b00010101000100011110: color_data = 12'b000001101111;
20'b00010101000100011111: color_data = 12'b000001101111;
20'b00010101000100100000: color_data = 12'b000001101111;
20'b00010101000100100001: color_data = 12'b000001101111;
20'b00010101000100100010: color_data = 12'b000001101111;
20'b00010101000100100011: color_data = 12'b000001101111;
20'b00010101000100100100: color_data = 12'b000001101111;
20'b00010101000100101101: color_data = 12'b000011111111;
20'b00010101000100101110: color_data = 12'b000011111111;
20'b00010101000100101111: color_data = 12'b000011111111;
20'b00010101000100110000: color_data = 12'b000011111111;
20'b00010101000100110001: color_data = 12'b000011111111;
20'b00010101000100110010: color_data = 12'b000011111111;
20'b00010101000100110011: color_data = 12'b000011111111;
20'b00010101000100110100: color_data = 12'b000011111111;
20'b00010101000100110101: color_data = 12'b000011111111;
20'b00010101000100110110: color_data = 12'b000011111111;
20'b00010101000100110111: color_data = 12'b000011111111;
20'b00010101000100111000: color_data = 12'b000011111111;
20'b00010101000100111001: color_data = 12'b000011111111;
20'b00010101000100111010: color_data = 12'b000011111111;
20'b00010101000100111011: color_data = 12'b000011111111;
20'b00010101000100111100: color_data = 12'b000011111111;
20'b00010101000100111101: color_data = 12'b000011111111;
20'b00010101000100111110: color_data = 12'b000011111111;
20'b00010101000100111111: color_data = 12'b000011111111;
20'b00010101000101000000: color_data = 12'b000011111111;
20'b00010101000101000001: color_data = 12'b000011111111;
20'b00010101000101000010: color_data = 12'b000011111111;
20'b00010101000101000011: color_data = 12'b000011111111;
20'b00010101000101000100: color_data = 12'b000011111111;
20'b00010101000101000101: color_data = 12'b000011111111;
20'b00010101000101000110: color_data = 12'b000011111111;
20'b00010101000101000111: color_data = 12'b000011111111;
20'b00010101000101001000: color_data = 12'b000011111111;
20'b00010101000101001001: color_data = 12'b000011111111;
20'b00010101000101001010: color_data = 12'b000011111111;
20'b00010101000101001011: color_data = 12'b000011111111;
20'b00010101000101001100: color_data = 12'b000011111111;
20'b00010101000101001101: color_data = 12'b000011111111;
20'b00010101000101001110: color_data = 12'b000011111111;
20'b00010101000101001111: color_data = 12'b000011111111;
20'b00010101000101010000: color_data = 12'b000011111111;
20'b00010101000101010001: color_data = 12'b000011111111;
20'b00010101000101010010: color_data = 12'b000011111111;
20'b00010101000101010011: color_data = 12'b000011111111;
20'b00010101000101010100: color_data = 12'b000011111111;
20'b00010101000101010101: color_data = 12'b000011111111;
20'b00010101000101011111: color_data = 12'b111101110000;
20'b00010101000101100000: color_data = 12'b111101110000;
20'b00010101000101100001: color_data = 12'b111101110000;
20'b00010101000101100010: color_data = 12'b111101110000;
20'b00010101000101100011: color_data = 12'b111101110000;
20'b00010101000101100100: color_data = 12'b111101110000;
20'b00010101000101100101: color_data = 12'b111101110000;
20'b00010101000101100110: color_data = 12'b111101110000;
20'b00010101000101100111: color_data = 12'b111101110000;
20'b00010101000101101000: color_data = 12'b111101110000;
20'b00010101000101101001: color_data = 12'b111101110000;
20'b00010101000101101010: color_data = 12'b111101110000;
20'b00010101000101101011: color_data = 12'b111101110000;
20'b00010101000101101100: color_data = 12'b111101110000;
20'b00010101000101101101: color_data = 12'b111101110000;
20'b00010101000101101110: color_data = 12'b111101110000;
20'b00010101000101101111: color_data = 12'b111101110000;
20'b00010101000101110000: color_data = 12'b111101110000;
20'b00010101000101110001: color_data = 12'b111101110000;
20'b00010101000101110010: color_data = 12'b111101110000;
20'b00010101000101110011: color_data = 12'b111101110000;
20'b00010101000101110100: color_data = 12'b111101110000;
20'b00010101000101110101: color_data = 12'b111101110000;
20'b00010101000101110110: color_data = 12'b111101110000;
20'b00010101000101110111: color_data = 12'b111101110000;
20'b00010101000101111000: color_data = 12'b111101110000;
20'b00010101000101111001: color_data = 12'b111101110000;
20'b00010101000101111010: color_data = 12'b111101110000;
20'b00010101000101111011: color_data = 12'b111101110000;
20'b00010101000101111100: color_data = 12'b111101110000;
20'b00010101000101111101: color_data = 12'b111101110000;
20'b00010101000101111110: color_data = 12'b111101110000;
20'b00010101000110000111: color_data = 12'b000011110000;
20'b00010101000110001000: color_data = 12'b000011110000;
20'b00010101000110001001: color_data = 12'b000011110000;
20'b00010101000110001010: color_data = 12'b000011110000;
20'b00010101000110001011: color_data = 12'b000011110000;
20'b00010101000110001100: color_data = 12'b000011110000;
20'b00010101000110001101: color_data = 12'b000011110000;
20'b00010101000110001110: color_data = 12'b000011110000;
20'b00010101000110001111: color_data = 12'b000011110000;
20'b00010101000110011000: color_data = 12'b111100001111;
20'b00010101000110011001: color_data = 12'b111100001111;
20'b00010101000110011010: color_data = 12'b111100001111;
20'b00010101000110011011: color_data = 12'b111100001111;
20'b00010101000110011100: color_data = 12'b111100001111;
20'b00010101000110011101: color_data = 12'b111100001111;
20'b00010101000110011110: color_data = 12'b111100001111;
20'b00010101000110011111: color_data = 12'b111100001111;
20'b00010101000110100000: color_data = 12'b111100001111;
20'b00010101000110100001: color_data = 12'b111100001111;
20'b00010101000110100010: color_data = 12'b111100001111;
20'b00010101000110100011: color_data = 12'b111100001111;
20'b00010101000110100100: color_data = 12'b111100001111;
20'b00010101000110100101: color_data = 12'b111100001111;
20'b00010101000110100110: color_data = 12'b111100001111;
20'b00010101000110100111: color_data = 12'b111100001111;
20'b00010101000110101000: color_data = 12'b111100001111;
20'b00010101000110101001: color_data = 12'b111100001111;
20'b00010101000110101010: color_data = 12'b111100001111;
20'b00010101000110101011: color_data = 12'b111100001111;
20'b00010101000110101100: color_data = 12'b111100001111;
20'b00010101000110101101: color_data = 12'b111100001111;
20'b00010101000110101110: color_data = 12'b111100001111;
20'b00010101000110101111: color_data = 12'b111100001111;
20'b00010101000110110000: color_data = 12'b111100001111;
20'b00010101000110110001: color_data = 12'b111100001111;
20'b00010101000110110010: color_data = 12'b111100001111;
20'b00010101000110110011: color_data = 12'b111100001111;
20'b00010101000110110100: color_data = 12'b111100001111;
20'b00010101000110110101: color_data = 12'b111100001111;
20'b00010101000110110110: color_data = 12'b111100001111;
20'b00010101000110110111: color_data = 12'b111100001111;
20'b00010101010011010011: color_data = 12'b000000001111;
20'b00010101010011010100: color_data = 12'b000000001111;
20'b00010101010011010101: color_data = 12'b000000001111;
20'b00010101010011010110: color_data = 12'b000000001111;
20'b00010101010011010111: color_data = 12'b000000001111;
20'b00010101010011011000: color_data = 12'b000000001111;
20'b00010101010011011001: color_data = 12'b000000001111;
20'b00010101010011011010: color_data = 12'b000000001111;
20'b00010101010011011011: color_data = 12'b000000001111;
20'b00010101010011011100: color_data = 12'b000000001111;
20'b00010101010011011101: color_data = 12'b000000001111;
20'b00010101010011011110: color_data = 12'b000000001111;
20'b00010101010011011111: color_data = 12'b000000001111;
20'b00010101010011100000: color_data = 12'b000000001111;
20'b00010101010011100001: color_data = 12'b000000001111;
20'b00010101010011100010: color_data = 12'b000000001111;
20'b00010101010011100011: color_data = 12'b000000001111;
20'b00010101010011100100: color_data = 12'b000000001111;
20'b00010101010011100101: color_data = 12'b000000001111;
20'b00010101010011100110: color_data = 12'b000000001111;
20'b00010101010011100111: color_data = 12'b000000001111;
20'b00010101010011101000: color_data = 12'b000000001111;
20'b00010101010011101001: color_data = 12'b000000001111;
20'b00010101010011101010: color_data = 12'b000000001111;
20'b00010101010011101011: color_data = 12'b000000001111;
20'b00010101010011101100: color_data = 12'b000000001111;
20'b00010101010011101101: color_data = 12'b000000001111;
20'b00010101010011101110: color_data = 12'b000000001111;
20'b00010101010011101111: color_data = 12'b000000001111;
20'b00010101010011110000: color_data = 12'b000000001111;
20'b00010101010011110001: color_data = 12'b000000001111;
20'b00010101010011110010: color_data = 12'b000000001111;
20'b00010101010011110011: color_data = 12'b000000001111;
20'b00010101010011110100: color_data = 12'b000000001111;
20'b00010101010011110101: color_data = 12'b000000001111;
20'b00010101010011110110: color_data = 12'b000000001111;
20'b00010101010011110111: color_data = 12'b000000001111;
20'b00010101010011111000: color_data = 12'b000000001111;
20'b00010101010011111001: color_data = 12'b000000001111;
20'b00010101010011111010: color_data = 12'b000000001111;
20'b00010101010011111011: color_data = 12'b000000001111;
20'b00010101010100000101: color_data = 12'b000001101111;
20'b00010101010100000110: color_data = 12'b000001101111;
20'b00010101010100000111: color_data = 12'b000001101111;
20'b00010101010100001000: color_data = 12'b000001101111;
20'b00010101010100001001: color_data = 12'b000001101111;
20'b00010101010100001010: color_data = 12'b000001101111;
20'b00010101010100001011: color_data = 12'b000001101111;
20'b00010101010100001100: color_data = 12'b000001101111;
20'b00010101010100001101: color_data = 12'b000001101111;
20'b00010101010100001110: color_data = 12'b000001101111;
20'b00010101010100001111: color_data = 12'b000001101111;
20'b00010101010100010000: color_data = 12'b000001101111;
20'b00010101010100010001: color_data = 12'b000001101111;
20'b00010101010100010010: color_data = 12'b000001101111;
20'b00010101010100010011: color_data = 12'b000001101111;
20'b00010101010100010100: color_data = 12'b000001101111;
20'b00010101010100010101: color_data = 12'b000001101111;
20'b00010101010100010110: color_data = 12'b000001101111;
20'b00010101010100010111: color_data = 12'b000001101111;
20'b00010101010100011000: color_data = 12'b000001101111;
20'b00010101010100011001: color_data = 12'b000001101111;
20'b00010101010100011010: color_data = 12'b000001101111;
20'b00010101010100011011: color_data = 12'b000001101111;
20'b00010101010100011100: color_data = 12'b000001101111;
20'b00010101010100011101: color_data = 12'b000001101111;
20'b00010101010100011110: color_data = 12'b000001101111;
20'b00010101010100011111: color_data = 12'b000001101111;
20'b00010101010100100000: color_data = 12'b000001101111;
20'b00010101010100100001: color_data = 12'b000001101111;
20'b00010101010100100010: color_data = 12'b000001101111;
20'b00010101010100100011: color_data = 12'b000001101111;
20'b00010101010100100100: color_data = 12'b000001101111;
20'b00010101010100101101: color_data = 12'b000011111111;
20'b00010101010100101110: color_data = 12'b000011111111;
20'b00010101010100101111: color_data = 12'b000011111111;
20'b00010101010100110000: color_data = 12'b000011111111;
20'b00010101010100110001: color_data = 12'b000011111111;
20'b00010101010100110010: color_data = 12'b000011111111;
20'b00010101010100110011: color_data = 12'b000011111111;
20'b00010101010100110100: color_data = 12'b000011111111;
20'b00010101010100110101: color_data = 12'b000011111111;
20'b00010101010100110110: color_data = 12'b000011111111;
20'b00010101010100110111: color_data = 12'b000011111111;
20'b00010101010100111000: color_data = 12'b000011111111;
20'b00010101010100111001: color_data = 12'b000011111111;
20'b00010101010100111010: color_data = 12'b000011111111;
20'b00010101010100111011: color_data = 12'b000011111111;
20'b00010101010100111100: color_data = 12'b000011111111;
20'b00010101010100111101: color_data = 12'b000011111111;
20'b00010101010100111110: color_data = 12'b000011111111;
20'b00010101010100111111: color_data = 12'b000011111111;
20'b00010101010101000000: color_data = 12'b000011111111;
20'b00010101010101000001: color_data = 12'b000011111111;
20'b00010101010101000010: color_data = 12'b000011111111;
20'b00010101010101000011: color_data = 12'b000011111111;
20'b00010101010101000100: color_data = 12'b000011111111;
20'b00010101010101000101: color_data = 12'b000011111111;
20'b00010101010101000110: color_data = 12'b000011111111;
20'b00010101010101000111: color_data = 12'b000011111111;
20'b00010101010101001000: color_data = 12'b000011111111;
20'b00010101010101001001: color_data = 12'b000011111111;
20'b00010101010101001010: color_data = 12'b000011111111;
20'b00010101010101001011: color_data = 12'b000011111111;
20'b00010101010101001100: color_data = 12'b000011111111;
20'b00010101010101001101: color_data = 12'b000011111111;
20'b00010101010101001110: color_data = 12'b000011111111;
20'b00010101010101001111: color_data = 12'b000011111111;
20'b00010101010101010000: color_data = 12'b000011111111;
20'b00010101010101010001: color_data = 12'b000011111111;
20'b00010101010101010010: color_data = 12'b000011111111;
20'b00010101010101010011: color_data = 12'b000011111111;
20'b00010101010101010100: color_data = 12'b000011111111;
20'b00010101010101010101: color_data = 12'b000011111111;
20'b00010101010101011111: color_data = 12'b111101110000;
20'b00010101010101100000: color_data = 12'b111101110000;
20'b00010101010101100001: color_data = 12'b111101110000;
20'b00010101010101100010: color_data = 12'b111101110000;
20'b00010101010101100011: color_data = 12'b111101110000;
20'b00010101010101100100: color_data = 12'b111101110000;
20'b00010101010101100101: color_data = 12'b111101110000;
20'b00010101010101100110: color_data = 12'b111101110000;
20'b00010101010101100111: color_data = 12'b111101110000;
20'b00010101010101101000: color_data = 12'b111101110000;
20'b00010101010101101001: color_data = 12'b111101110000;
20'b00010101010101101010: color_data = 12'b111101110000;
20'b00010101010101101011: color_data = 12'b111101110000;
20'b00010101010101101100: color_data = 12'b111101110000;
20'b00010101010101101101: color_data = 12'b111101110000;
20'b00010101010101101110: color_data = 12'b111101110000;
20'b00010101010101101111: color_data = 12'b111101110000;
20'b00010101010101110000: color_data = 12'b111101110000;
20'b00010101010101110001: color_data = 12'b111101110000;
20'b00010101010101110010: color_data = 12'b111101110000;
20'b00010101010101110011: color_data = 12'b111101110000;
20'b00010101010101110100: color_data = 12'b111101110000;
20'b00010101010101110101: color_data = 12'b111101110000;
20'b00010101010101110110: color_data = 12'b111101110000;
20'b00010101010101110111: color_data = 12'b111101110000;
20'b00010101010101111000: color_data = 12'b111101110000;
20'b00010101010101111001: color_data = 12'b111101110000;
20'b00010101010101111010: color_data = 12'b111101110000;
20'b00010101010101111011: color_data = 12'b111101110000;
20'b00010101010101111100: color_data = 12'b111101110000;
20'b00010101010101111101: color_data = 12'b111101110000;
20'b00010101010101111110: color_data = 12'b111101110000;
20'b00010101010110000111: color_data = 12'b000011110000;
20'b00010101010110001000: color_data = 12'b000011110000;
20'b00010101010110001001: color_data = 12'b000011110000;
20'b00010101010110001010: color_data = 12'b000011110000;
20'b00010101010110001011: color_data = 12'b000011110000;
20'b00010101010110001100: color_data = 12'b000011110000;
20'b00010101010110001101: color_data = 12'b000011110000;
20'b00010101010110001110: color_data = 12'b000011110000;
20'b00010101010110001111: color_data = 12'b000011110000;
20'b00010101010110011000: color_data = 12'b111100001111;
20'b00010101010110011001: color_data = 12'b111100001111;
20'b00010101010110011010: color_data = 12'b111100001111;
20'b00010101010110011011: color_data = 12'b111100001111;
20'b00010101010110011100: color_data = 12'b111100001111;
20'b00010101010110011101: color_data = 12'b111100001111;
20'b00010101010110011110: color_data = 12'b111100001111;
20'b00010101010110011111: color_data = 12'b111100001111;
20'b00010101010110100000: color_data = 12'b111100001111;
20'b00010101010110100001: color_data = 12'b111100001111;
20'b00010101010110100010: color_data = 12'b111100001111;
20'b00010101010110100011: color_data = 12'b111100001111;
20'b00010101010110100100: color_data = 12'b111100001111;
20'b00010101010110100101: color_data = 12'b111100001111;
20'b00010101010110100110: color_data = 12'b111100001111;
20'b00010101010110100111: color_data = 12'b111100001111;
20'b00010101010110101000: color_data = 12'b111100001111;
20'b00010101010110101001: color_data = 12'b111100001111;
20'b00010101010110101010: color_data = 12'b111100001111;
20'b00010101010110101011: color_data = 12'b111100001111;
20'b00010101010110101100: color_data = 12'b111100001111;
20'b00010101010110101101: color_data = 12'b111100001111;
20'b00010101010110101110: color_data = 12'b111100001111;
20'b00010101010110101111: color_data = 12'b111100001111;
20'b00010101010110110000: color_data = 12'b111100001111;
20'b00010101010110110001: color_data = 12'b111100001111;
20'b00010101010110110010: color_data = 12'b111100001111;
20'b00010101010110110011: color_data = 12'b111100001111;
20'b00010101010110110100: color_data = 12'b111100001111;
20'b00010101010110110101: color_data = 12'b111100001111;
20'b00010101010110110110: color_data = 12'b111100001111;
20'b00010101010110110111: color_data = 12'b111100001111;
20'b00010101100011010011: color_data = 12'b000000001111;
20'b00010101100011010100: color_data = 12'b000000001111;
20'b00010101100011010101: color_data = 12'b000000001111;
20'b00010101100011010110: color_data = 12'b000000001111;
20'b00010101100011010111: color_data = 12'b000000001111;
20'b00010101100011011000: color_data = 12'b000000001111;
20'b00010101100011011001: color_data = 12'b000000001111;
20'b00010101100011011010: color_data = 12'b000000001111;
20'b00010101100011011011: color_data = 12'b000000001111;
20'b00010101100011011100: color_data = 12'b000000001111;
20'b00010101100011011101: color_data = 12'b000000001111;
20'b00010101100011011110: color_data = 12'b000000001111;
20'b00010101100011011111: color_data = 12'b000000001111;
20'b00010101100011100000: color_data = 12'b000000001111;
20'b00010101100011100001: color_data = 12'b000000001111;
20'b00010101100011100010: color_data = 12'b000000001111;
20'b00010101100011100011: color_data = 12'b000000001111;
20'b00010101100011100100: color_data = 12'b000000001111;
20'b00010101100011100101: color_data = 12'b000000001111;
20'b00010101100011100110: color_data = 12'b000000001111;
20'b00010101100011100111: color_data = 12'b000000001111;
20'b00010101100011101000: color_data = 12'b000000001111;
20'b00010101100011101001: color_data = 12'b000000001111;
20'b00010101100011101010: color_data = 12'b000000001111;
20'b00010101100011101011: color_data = 12'b000000001111;
20'b00010101100011101100: color_data = 12'b000000001111;
20'b00010101100011101101: color_data = 12'b000000001111;
20'b00010101100011101110: color_data = 12'b000000001111;
20'b00010101100011101111: color_data = 12'b000000001111;
20'b00010101100011110000: color_data = 12'b000000001111;
20'b00010101100011110001: color_data = 12'b000000001111;
20'b00010101100011110010: color_data = 12'b000000001111;
20'b00010101100011110011: color_data = 12'b000000001111;
20'b00010101100011110100: color_data = 12'b000000001111;
20'b00010101100011110101: color_data = 12'b000000001111;
20'b00010101100011110110: color_data = 12'b000000001111;
20'b00010101100011110111: color_data = 12'b000000001111;
20'b00010101100011111000: color_data = 12'b000000001111;
20'b00010101100011111001: color_data = 12'b000000001111;
20'b00010101100011111010: color_data = 12'b000000001111;
20'b00010101100011111011: color_data = 12'b000000001111;
20'b00010101100100000101: color_data = 12'b000001101111;
20'b00010101100100000110: color_data = 12'b000001101111;
20'b00010101100100000111: color_data = 12'b000001101111;
20'b00010101100100001000: color_data = 12'b000001101111;
20'b00010101100100001001: color_data = 12'b000001101111;
20'b00010101100100001010: color_data = 12'b000001101111;
20'b00010101100100001011: color_data = 12'b000001101111;
20'b00010101100100001100: color_data = 12'b000001101111;
20'b00010101100100001101: color_data = 12'b000001101111;
20'b00010101100100001110: color_data = 12'b000001101111;
20'b00010101100100001111: color_data = 12'b000001101111;
20'b00010101100100010000: color_data = 12'b000001101111;
20'b00010101100100010001: color_data = 12'b000001101111;
20'b00010101100100010010: color_data = 12'b000001101111;
20'b00010101100100010011: color_data = 12'b000001101111;
20'b00010101100100010100: color_data = 12'b000001101111;
20'b00010101100100010101: color_data = 12'b000001101111;
20'b00010101100100010110: color_data = 12'b000001101111;
20'b00010101100100010111: color_data = 12'b000001101111;
20'b00010101100100011000: color_data = 12'b000001101111;
20'b00010101100100011001: color_data = 12'b000001101111;
20'b00010101100100011010: color_data = 12'b000001101111;
20'b00010101100100011011: color_data = 12'b000001101111;
20'b00010101100100011100: color_data = 12'b000001101111;
20'b00010101100100011101: color_data = 12'b000001101111;
20'b00010101100100011110: color_data = 12'b000001101111;
20'b00010101100100011111: color_data = 12'b000001101111;
20'b00010101100100100000: color_data = 12'b000001101111;
20'b00010101100100100001: color_data = 12'b000001101111;
20'b00010101100100100010: color_data = 12'b000001101111;
20'b00010101100100100011: color_data = 12'b000001101111;
20'b00010101100100100100: color_data = 12'b000001101111;
20'b00010101100100101101: color_data = 12'b000011111111;
20'b00010101100100101110: color_data = 12'b000011111111;
20'b00010101100100101111: color_data = 12'b000011111111;
20'b00010101100100110000: color_data = 12'b000011111111;
20'b00010101100100110001: color_data = 12'b000011111111;
20'b00010101100100110010: color_data = 12'b000011111111;
20'b00010101100100110011: color_data = 12'b000011111111;
20'b00010101100100110100: color_data = 12'b000011111111;
20'b00010101100100110101: color_data = 12'b000011111111;
20'b00010101100100110110: color_data = 12'b000011111111;
20'b00010101100100110111: color_data = 12'b000011111111;
20'b00010101100100111000: color_data = 12'b000011111111;
20'b00010101100100111001: color_data = 12'b000011111111;
20'b00010101100100111010: color_data = 12'b000011111111;
20'b00010101100100111011: color_data = 12'b000011111111;
20'b00010101100100111100: color_data = 12'b000011111111;
20'b00010101100100111101: color_data = 12'b000011111111;
20'b00010101100100111110: color_data = 12'b000011111111;
20'b00010101100100111111: color_data = 12'b000011111111;
20'b00010101100101000000: color_data = 12'b000011111111;
20'b00010101100101000001: color_data = 12'b000011111111;
20'b00010101100101000010: color_data = 12'b000011111111;
20'b00010101100101000011: color_data = 12'b000011111111;
20'b00010101100101000100: color_data = 12'b000011111111;
20'b00010101100101000101: color_data = 12'b000011111111;
20'b00010101100101000110: color_data = 12'b000011111111;
20'b00010101100101000111: color_data = 12'b000011111111;
20'b00010101100101001000: color_data = 12'b000011111111;
20'b00010101100101001001: color_data = 12'b000011111111;
20'b00010101100101001010: color_data = 12'b000011111111;
20'b00010101100101001011: color_data = 12'b000011111111;
20'b00010101100101001100: color_data = 12'b000011111111;
20'b00010101100101001101: color_data = 12'b000011111111;
20'b00010101100101001110: color_data = 12'b000011111111;
20'b00010101100101001111: color_data = 12'b000011111111;
20'b00010101100101010000: color_data = 12'b000011111111;
20'b00010101100101010001: color_data = 12'b000011111111;
20'b00010101100101010010: color_data = 12'b000011111111;
20'b00010101100101010011: color_data = 12'b000011111111;
20'b00010101100101010100: color_data = 12'b000011111111;
20'b00010101100101010101: color_data = 12'b000011111111;
20'b00010101100101011111: color_data = 12'b111101110000;
20'b00010101100101100000: color_data = 12'b111101110000;
20'b00010101100101100001: color_data = 12'b111101110000;
20'b00010101100101100010: color_data = 12'b111101110000;
20'b00010101100101100011: color_data = 12'b111101110000;
20'b00010101100101100100: color_data = 12'b111101110000;
20'b00010101100101100101: color_data = 12'b111101110000;
20'b00010101100101100110: color_data = 12'b111101110000;
20'b00010101100101100111: color_data = 12'b111101110000;
20'b00010101100101101000: color_data = 12'b111101110000;
20'b00010101100101101001: color_data = 12'b111101110000;
20'b00010101100101101010: color_data = 12'b111101110000;
20'b00010101100101101011: color_data = 12'b111101110000;
20'b00010101100101101100: color_data = 12'b111101110000;
20'b00010101100101101101: color_data = 12'b111101110000;
20'b00010101100101101110: color_data = 12'b111101110000;
20'b00010101100101101111: color_data = 12'b111101110000;
20'b00010101100101110000: color_data = 12'b111101110000;
20'b00010101100101110001: color_data = 12'b111101110000;
20'b00010101100101110010: color_data = 12'b111101110000;
20'b00010101100101110011: color_data = 12'b111101110000;
20'b00010101100101110100: color_data = 12'b111101110000;
20'b00010101100101110101: color_data = 12'b111101110000;
20'b00010101100101110110: color_data = 12'b111101110000;
20'b00010101100101110111: color_data = 12'b111101110000;
20'b00010101100101111000: color_data = 12'b111101110000;
20'b00010101100101111001: color_data = 12'b111101110000;
20'b00010101100101111010: color_data = 12'b111101110000;
20'b00010101100101111011: color_data = 12'b111101110000;
20'b00010101100101111100: color_data = 12'b111101110000;
20'b00010101100101111101: color_data = 12'b111101110000;
20'b00010101100101111110: color_data = 12'b111101110000;
20'b00010101100110000111: color_data = 12'b000011110000;
20'b00010101100110001000: color_data = 12'b000011110000;
20'b00010101100110001001: color_data = 12'b000011110000;
20'b00010101100110001010: color_data = 12'b000011110000;
20'b00010101100110001011: color_data = 12'b000011110000;
20'b00010101100110001100: color_data = 12'b000011110000;
20'b00010101100110001101: color_data = 12'b000011110000;
20'b00010101100110001110: color_data = 12'b000011110000;
20'b00010101100110001111: color_data = 12'b000011110000;
20'b00010101100110011000: color_data = 12'b111100001111;
20'b00010101100110011001: color_data = 12'b111100001111;
20'b00010101100110011010: color_data = 12'b111100001111;
20'b00010101100110011011: color_data = 12'b111100001111;
20'b00010101100110011100: color_data = 12'b111100001111;
20'b00010101100110011101: color_data = 12'b111100001111;
20'b00010101100110011110: color_data = 12'b111100001111;
20'b00010101100110011111: color_data = 12'b111100001111;
20'b00010101100110100000: color_data = 12'b111100001111;
20'b00010101100110100001: color_data = 12'b111100001111;
20'b00010101100110100010: color_data = 12'b111100001111;
20'b00010101100110100011: color_data = 12'b111100001111;
20'b00010101100110100100: color_data = 12'b111100001111;
20'b00010101100110100101: color_data = 12'b111100001111;
20'b00010101100110100110: color_data = 12'b111100001111;
20'b00010101100110100111: color_data = 12'b111100001111;
20'b00010101100110101000: color_data = 12'b111100001111;
20'b00010101100110101001: color_data = 12'b111100001111;
20'b00010101100110101010: color_data = 12'b111100001111;
20'b00010101100110101011: color_data = 12'b111100001111;
20'b00010101100110101100: color_data = 12'b111100001111;
20'b00010101100110101101: color_data = 12'b111100001111;
20'b00010101100110101110: color_data = 12'b111100001111;
20'b00010101100110101111: color_data = 12'b111100001111;
20'b00010101100110110000: color_data = 12'b111100001111;
20'b00010101100110110001: color_data = 12'b111100001111;
20'b00010101100110110010: color_data = 12'b111100001111;
20'b00010101100110110011: color_data = 12'b111100001111;
20'b00010101100110110100: color_data = 12'b111100001111;
20'b00010101100110110101: color_data = 12'b111100001111;
20'b00010101100110110110: color_data = 12'b111100001111;
20'b00010101100110110111: color_data = 12'b111100001111;
20'b00010101110011010011: color_data = 12'b000000001111;
20'b00010101110011010100: color_data = 12'b000000001111;
20'b00010101110011010101: color_data = 12'b000000001111;
20'b00010101110011010110: color_data = 12'b000000001111;
20'b00010101110011010111: color_data = 12'b000000001111;
20'b00010101110011011000: color_data = 12'b000000001111;
20'b00010101110011011001: color_data = 12'b000000001111;
20'b00010101110011011010: color_data = 12'b000000001111;
20'b00010101110011011011: color_data = 12'b000000001111;
20'b00010101110011011100: color_data = 12'b000000001111;
20'b00010101110011011101: color_data = 12'b000000001111;
20'b00010101110011011110: color_data = 12'b000000001111;
20'b00010101110011011111: color_data = 12'b000000001111;
20'b00010101110011100000: color_data = 12'b000000001111;
20'b00010101110011100001: color_data = 12'b000000001111;
20'b00010101110011100010: color_data = 12'b000000001111;
20'b00010101110011100011: color_data = 12'b000000001111;
20'b00010101110011100100: color_data = 12'b000000001111;
20'b00010101110011100101: color_data = 12'b000000001111;
20'b00010101110011100110: color_data = 12'b000000001111;
20'b00010101110011100111: color_data = 12'b000000001111;
20'b00010101110011101000: color_data = 12'b000000001111;
20'b00010101110011101001: color_data = 12'b000000001111;
20'b00010101110011101010: color_data = 12'b000000001111;
20'b00010101110011101011: color_data = 12'b000000001111;
20'b00010101110011101100: color_data = 12'b000000001111;
20'b00010101110011101101: color_data = 12'b000000001111;
20'b00010101110011101110: color_data = 12'b000000001111;
20'b00010101110011101111: color_data = 12'b000000001111;
20'b00010101110011110000: color_data = 12'b000000001111;
20'b00010101110011110001: color_data = 12'b000000001111;
20'b00010101110011110010: color_data = 12'b000000001111;
20'b00010101110011110011: color_data = 12'b000000001111;
20'b00010101110011110100: color_data = 12'b000000001111;
20'b00010101110011110101: color_data = 12'b000000001111;
20'b00010101110011110110: color_data = 12'b000000001111;
20'b00010101110011110111: color_data = 12'b000000001111;
20'b00010101110011111000: color_data = 12'b000000001111;
20'b00010101110011111001: color_data = 12'b000000001111;
20'b00010101110011111010: color_data = 12'b000000001111;
20'b00010101110011111011: color_data = 12'b000000001111;
20'b00010101110100000101: color_data = 12'b000001101111;
20'b00010101110100000110: color_data = 12'b000001101111;
20'b00010101110100000111: color_data = 12'b000001101111;
20'b00010101110100001000: color_data = 12'b000001101111;
20'b00010101110100001001: color_data = 12'b000001101111;
20'b00010101110100001010: color_data = 12'b000001101111;
20'b00010101110100001011: color_data = 12'b000001101111;
20'b00010101110100001100: color_data = 12'b000001101111;
20'b00010101110100001101: color_data = 12'b000001101111;
20'b00010101110100001110: color_data = 12'b000001101111;
20'b00010101110100001111: color_data = 12'b000001101111;
20'b00010101110100010000: color_data = 12'b000001101111;
20'b00010101110100010001: color_data = 12'b000001101111;
20'b00010101110100010010: color_data = 12'b000001101111;
20'b00010101110100010011: color_data = 12'b000001101111;
20'b00010101110100010100: color_data = 12'b000001101111;
20'b00010101110100010101: color_data = 12'b000001101111;
20'b00010101110100010110: color_data = 12'b000001101111;
20'b00010101110100010111: color_data = 12'b000001101111;
20'b00010101110100011000: color_data = 12'b000001101111;
20'b00010101110100011001: color_data = 12'b000001101111;
20'b00010101110100011010: color_data = 12'b000001101111;
20'b00010101110100011011: color_data = 12'b000001101111;
20'b00010101110100011100: color_data = 12'b000001101111;
20'b00010101110100011101: color_data = 12'b000001101111;
20'b00010101110100011110: color_data = 12'b000001101111;
20'b00010101110100011111: color_data = 12'b000001101111;
20'b00010101110100100000: color_data = 12'b000001101111;
20'b00010101110100100001: color_data = 12'b000001101111;
20'b00010101110100100010: color_data = 12'b000001101111;
20'b00010101110100100011: color_data = 12'b000001101111;
20'b00010101110100100100: color_data = 12'b000001101111;
20'b00010101110100101101: color_data = 12'b000011111111;
20'b00010101110100101110: color_data = 12'b000011111111;
20'b00010101110100101111: color_data = 12'b000011111111;
20'b00010101110100110000: color_data = 12'b000011111111;
20'b00010101110100110001: color_data = 12'b000011111111;
20'b00010101110100110010: color_data = 12'b000011111111;
20'b00010101110100110011: color_data = 12'b000011111111;
20'b00010101110100110100: color_data = 12'b000011111111;
20'b00010101110100110101: color_data = 12'b000011111111;
20'b00010101110100110110: color_data = 12'b000011111111;
20'b00010101110100110111: color_data = 12'b000011111111;
20'b00010101110100111000: color_data = 12'b000011111111;
20'b00010101110100111001: color_data = 12'b000011111111;
20'b00010101110100111010: color_data = 12'b000011111111;
20'b00010101110100111011: color_data = 12'b000011111111;
20'b00010101110100111100: color_data = 12'b000011111111;
20'b00010101110100111101: color_data = 12'b000011111111;
20'b00010101110100111110: color_data = 12'b000011111111;
20'b00010101110100111111: color_data = 12'b000011111111;
20'b00010101110101000000: color_data = 12'b000011111111;
20'b00010101110101000001: color_data = 12'b000011111111;
20'b00010101110101000010: color_data = 12'b000011111111;
20'b00010101110101000011: color_data = 12'b000011111111;
20'b00010101110101000100: color_data = 12'b000011111111;
20'b00010101110101000101: color_data = 12'b000011111111;
20'b00010101110101000110: color_data = 12'b000011111111;
20'b00010101110101000111: color_data = 12'b000011111111;
20'b00010101110101001000: color_data = 12'b000011111111;
20'b00010101110101001001: color_data = 12'b000011111111;
20'b00010101110101001010: color_data = 12'b000011111111;
20'b00010101110101001011: color_data = 12'b000011111111;
20'b00010101110101001100: color_data = 12'b000011111111;
20'b00010101110101001101: color_data = 12'b000011111111;
20'b00010101110101001110: color_data = 12'b000011111111;
20'b00010101110101001111: color_data = 12'b000011111111;
20'b00010101110101010000: color_data = 12'b000011111111;
20'b00010101110101010001: color_data = 12'b000011111111;
20'b00010101110101010010: color_data = 12'b000011111111;
20'b00010101110101010011: color_data = 12'b000011111111;
20'b00010101110101010100: color_data = 12'b000011111111;
20'b00010101110101010101: color_data = 12'b000011111111;
20'b00010101110101011111: color_data = 12'b111101110000;
20'b00010101110101100000: color_data = 12'b111101110000;
20'b00010101110101100001: color_data = 12'b111101110000;
20'b00010101110101100010: color_data = 12'b111101110000;
20'b00010101110101100011: color_data = 12'b111101110000;
20'b00010101110101100100: color_data = 12'b111101110000;
20'b00010101110101100101: color_data = 12'b111101110000;
20'b00010101110101100110: color_data = 12'b111101110000;
20'b00010101110101100111: color_data = 12'b111101110000;
20'b00010101110101101000: color_data = 12'b111101110000;
20'b00010101110101101001: color_data = 12'b111101110000;
20'b00010101110101101010: color_data = 12'b111101110000;
20'b00010101110101101011: color_data = 12'b111101110000;
20'b00010101110101101100: color_data = 12'b111101110000;
20'b00010101110101101101: color_data = 12'b111101110000;
20'b00010101110101101110: color_data = 12'b111101110000;
20'b00010101110101101111: color_data = 12'b111101110000;
20'b00010101110101110000: color_data = 12'b111101110000;
20'b00010101110101110001: color_data = 12'b111101110000;
20'b00010101110101110010: color_data = 12'b111101110000;
20'b00010101110101110011: color_data = 12'b111101110000;
20'b00010101110101110100: color_data = 12'b111101110000;
20'b00010101110101110101: color_data = 12'b111101110000;
20'b00010101110101110110: color_data = 12'b111101110000;
20'b00010101110101110111: color_data = 12'b111101110000;
20'b00010101110101111000: color_data = 12'b111101110000;
20'b00010101110101111001: color_data = 12'b111101110000;
20'b00010101110101111010: color_data = 12'b111101110000;
20'b00010101110101111011: color_data = 12'b111101110000;
20'b00010101110101111100: color_data = 12'b111101110000;
20'b00010101110101111101: color_data = 12'b111101110000;
20'b00010101110101111110: color_data = 12'b111101110000;
20'b00010101110110000111: color_data = 12'b000011110000;
20'b00010101110110001000: color_data = 12'b000011110000;
20'b00010101110110001001: color_data = 12'b000011110000;
20'b00010101110110001010: color_data = 12'b000011110000;
20'b00010101110110001011: color_data = 12'b000011110000;
20'b00010101110110001100: color_data = 12'b000011110000;
20'b00010101110110001101: color_data = 12'b000011110000;
20'b00010101110110001110: color_data = 12'b000011110000;
20'b00010101110110001111: color_data = 12'b000011110000;
20'b00010101110110011000: color_data = 12'b111100001111;
20'b00010101110110011001: color_data = 12'b111100001111;
20'b00010101110110011010: color_data = 12'b111100001111;
20'b00010101110110011011: color_data = 12'b111100001111;
20'b00010101110110011100: color_data = 12'b111100001111;
20'b00010101110110011101: color_data = 12'b111100001111;
20'b00010101110110011110: color_data = 12'b111100001111;
20'b00010101110110011111: color_data = 12'b111100001111;
20'b00010101110110100000: color_data = 12'b111100001111;
20'b00010101110110100001: color_data = 12'b111100001111;
20'b00010101110110100010: color_data = 12'b111100001111;
20'b00010101110110100011: color_data = 12'b111100001111;
20'b00010101110110100100: color_data = 12'b111100001111;
20'b00010101110110100101: color_data = 12'b111100001111;
20'b00010101110110100110: color_data = 12'b111100001111;
20'b00010101110110100111: color_data = 12'b111100001111;
20'b00010101110110101000: color_data = 12'b111100001111;
20'b00010101110110101001: color_data = 12'b111100001111;
20'b00010101110110101010: color_data = 12'b111100001111;
20'b00010101110110101011: color_data = 12'b111100001111;
20'b00010101110110101100: color_data = 12'b111100001111;
20'b00010101110110101101: color_data = 12'b111100001111;
20'b00010101110110101110: color_data = 12'b111100001111;
20'b00010101110110101111: color_data = 12'b111100001111;
20'b00010101110110110000: color_data = 12'b111100001111;
20'b00010101110110110001: color_data = 12'b111100001111;
20'b00010101110110110010: color_data = 12'b111100001111;
20'b00010101110110110011: color_data = 12'b111100001111;
20'b00010101110110110100: color_data = 12'b111100001111;
20'b00010101110110110101: color_data = 12'b111100001111;
20'b00010101110110110110: color_data = 12'b111100001111;
20'b00010101110110110111: color_data = 12'b111100001111;
20'b00010110000011010011: color_data = 12'b000000001111;
20'b00010110000011010100: color_data = 12'b000000001111;
20'b00010110000011010101: color_data = 12'b000000001111;
20'b00010110000011010110: color_data = 12'b000000001111;
20'b00010110000011010111: color_data = 12'b000000001111;
20'b00010110000011011000: color_data = 12'b000000001111;
20'b00010110000011011001: color_data = 12'b000000001111;
20'b00010110000011011010: color_data = 12'b000000001111;
20'b00010110000011011011: color_data = 12'b000000001111;
20'b00010110000011011100: color_data = 12'b000000001111;
20'b00010110000011011101: color_data = 12'b000000001111;
20'b00010110000011011110: color_data = 12'b000000001111;
20'b00010110000011011111: color_data = 12'b000000001111;
20'b00010110000011100000: color_data = 12'b000000001111;
20'b00010110000011100001: color_data = 12'b000000001111;
20'b00010110000011100010: color_data = 12'b000000001111;
20'b00010110000011100011: color_data = 12'b000000001111;
20'b00010110000011100100: color_data = 12'b000000001111;
20'b00010110000011100101: color_data = 12'b000000001111;
20'b00010110000011100110: color_data = 12'b000000001111;
20'b00010110000011100111: color_data = 12'b000000001111;
20'b00010110000011101000: color_data = 12'b000000001111;
20'b00010110000011101001: color_data = 12'b000000001111;
20'b00010110000011101010: color_data = 12'b000000001111;
20'b00010110000011101011: color_data = 12'b000000001111;
20'b00010110000011101100: color_data = 12'b000000001111;
20'b00010110000011101101: color_data = 12'b000000001111;
20'b00010110000011101110: color_data = 12'b000000001111;
20'b00010110000011101111: color_data = 12'b000000001111;
20'b00010110000011110000: color_data = 12'b000000001111;
20'b00010110000011110001: color_data = 12'b000000001111;
20'b00010110000011110010: color_data = 12'b000000001111;
20'b00010110000011110011: color_data = 12'b000000001111;
20'b00010110000011110100: color_data = 12'b000000001111;
20'b00010110000011110101: color_data = 12'b000000001111;
20'b00010110000011110110: color_data = 12'b000000001111;
20'b00010110000011110111: color_data = 12'b000000001111;
20'b00010110000011111000: color_data = 12'b000000001111;
20'b00010110000011111001: color_data = 12'b000000001111;
20'b00010110000011111010: color_data = 12'b000000001111;
20'b00010110000011111011: color_data = 12'b000000001111;
20'b00010110000100000101: color_data = 12'b000001101111;
20'b00010110000100000110: color_data = 12'b000001101111;
20'b00010110000100000111: color_data = 12'b000001101111;
20'b00010110000100001000: color_data = 12'b000001101111;
20'b00010110000100001001: color_data = 12'b000001101111;
20'b00010110000100001010: color_data = 12'b000001101111;
20'b00010110000100001011: color_data = 12'b000001101111;
20'b00010110000100001100: color_data = 12'b000001101111;
20'b00010110000100001101: color_data = 12'b000001101111;
20'b00010110000100001110: color_data = 12'b000001101111;
20'b00010110000100001111: color_data = 12'b000001101111;
20'b00010110000100010000: color_data = 12'b000001101111;
20'b00010110000100010001: color_data = 12'b000001101111;
20'b00010110000100010010: color_data = 12'b000001101111;
20'b00010110000100010011: color_data = 12'b000001101111;
20'b00010110000100010100: color_data = 12'b000001101111;
20'b00010110000100010101: color_data = 12'b000001101111;
20'b00010110000100010110: color_data = 12'b000001101111;
20'b00010110000100010111: color_data = 12'b000001101111;
20'b00010110000100011000: color_data = 12'b000001101111;
20'b00010110000100011001: color_data = 12'b000001101111;
20'b00010110000100011010: color_data = 12'b000001101111;
20'b00010110000100011011: color_data = 12'b000001101111;
20'b00010110000100011100: color_data = 12'b000001101111;
20'b00010110000100011101: color_data = 12'b000001101111;
20'b00010110000100011110: color_data = 12'b000001101111;
20'b00010110000100011111: color_data = 12'b000001101111;
20'b00010110000100100000: color_data = 12'b000001101111;
20'b00010110000100100001: color_data = 12'b000001101111;
20'b00010110000100100010: color_data = 12'b000001101111;
20'b00010110000100100011: color_data = 12'b000001101111;
20'b00010110000100100100: color_data = 12'b000001101111;
20'b00010110000100101101: color_data = 12'b000011111111;
20'b00010110000100101110: color_data = 12'b000011111111;
20'b00010110000100101111: color_data = 12'b000011111111;
20'b00010110000100110000: color_data = 12'b000011111111;
20'b00010110000100110001: color_data = 12'b000011111111;
20'b00010110000100110010: color_data = 12'b000011111111;
20'b00010110000100110011: color_data = 12'b000011111111;
20'b00010110000100110100: color_data = 12'b000011111111;
20'b00010110000100110101: color_data = 12'b000011111111;
20'b00010110000100110110: color_data = 12'b000011111111;
20'b00010110000100110111: color_data = 12'b000011111111;
20'b00010110000100111000: color_data = 12'b000011111111;
20'b00010110000100111001: color_data = 12'b000011111111;
20'b00010110000100111010: color_data = 12'b000011111111;
20'b00010110000100111011: color_data = 12'b000011111111;
20'b00010110000100111100: color_data = 12'b000011111111;
20'b00010110000100111101: color_data = 12'b000011111111;
20'b00010110000100111110: color_data = 12'b000011111111;
20'b00010110000100111111: color_data = 12'b000011111111;
20'b00010110000101000000: color_data = 12'b000011111111;
20'b00010110000101000001: color_data = 12'b000011111111;
20'b00010110000101000010: color_data = 12'b000011111111;
20'b00010110000101000011: color_data = 12'b000011111111;
20'b00010110000101000100: color_data = 12'b000011111111;
20'b00010110000101000101: color_data = 12'b000011111111;
20'b00010110000101000110: color_data = 12'b000011111111;
20'b00010110000101000111: color_data = 12'b000011111111;
20'b00010110000101001000: color_data = 12'b000011111111;
20'b00010110000101001001: color_data = 12'b000011111111;
20'b00010110000101001010: color_data = 12'b000011111111;
20'b00010110000101001011: color_data = 12'b000011111111;
20'b00010110000101001100: color_data = 12'b000011111111;
20'b00010110000101001101: color_data = 12'b000011111111;
20'b00010110000101001110: color_data = 12'b000011111111;
20'b00010110000101001111: color_data = 12'b000011111111;
20'b00010110000101010000: color_data = 12'b000011111111;
20'b00010110000101010001: color_data = 12'b000011111111;
20'b00010110000101010010: color_data = 12'b000011111111;
20'b00010110000101010011: color_data = 12'b000011111111;
20'b00010110000101010100: color_data = 12'b000011111111;
20'b00010110000101010101: color_data = 12'b000011111111;
20'b00010110000101011111: color_data = 12'b111101110000;
20'b00010110000101100000: color_data = 12'b111101110000;
20'b00010110000101100001: color_data = 12'b111101110000;
20'b00010110000101100010: color_data = 12'b111101110000;
20'b00010110000101100011: color_data = 12'b111101110000;
20'b00010110000101100100: color_data = 12'b111101110000;
20'b00010110000101100101: color_data = 12'b111101110000;
20'b00010110000101100110: color_data = 12'b111101110000;
20'b00010110000101100111: color_data = 12'b111101110000;
20'b00010110000101101000: color_data = 12'b111101110000;
20'b00010110000101101001: color_data = 12'b111101110000;
20'b00010110000101101010: color_data = 12'b111101110000;
20'b00010110000101101011: color_data = 12'b111101110000;
20'b00010110000101101100: color_data = 12'b111101110000;
20'b00010110000101101101: color_data = 12'b111101110000;
20'b00010110000101101110: color_data = 12'b111101110000;
20'b00010110000101101111: color_data = 12'b111101110000;
20'b00010110000101110000: color_data = 12'b111101110000;
20'b00010110000101110001: color_data = 12'b111101110000;
20'b00010110000101110010: color_data = 12'b111101110000;
20'b00010110000101110011: color_data = 12'b111101110000;
20'b00010110000101110100: color_data = 12'b111101110000;
20'b00010110000101110101: color_data = 12'b111101110000;
20'b00010110000101110110: color_data = 12'b111101110000;
20'b00010110000101110111: color_data = 12'b111101110000;
20'b00010110000101111000: color_data = 12'b111101110000;
20'b00010110000101111001: color_data = 12'b111101110000;
20'b00010110000101111010: color_data = 12'b111101110000;
20'b00010110000101111011: color_data = 12'b111101110000;
20'b00010110000101111100: color_data = 12'b111101110000;
20'b00010110000101111101: color_data = 12'b111101110000;
20'b00010110000101111110: color_data = 12'b111101110000;
20'b00010110000110000111: color_data = 12'b000011110000;
20'b00010110000110001000: color_data = 12'b000011110000;
20'b00010110000110001001: color_data = 12'b000011110000;
20'b00010110000110001010: color_data = 12'b000011110000;
20'b00010110000110001011: color_data = 12'b000011110000;
20'b00010110000110001100: color_data = 12'b000011110000;
20'b00010110000110001101: color_data = 12'b000011110000;
20'b00010110000110001110: color_data = 12'b000011110000;
20'b00010110000110001111: color_data = 12'b000011110000;
20'b00010110000110011000: color_data = 12'b111100001111;
20'b00010110000110011001: color_data = 12'b111100001111;
20'b00010110000110011010: color_data = 12'b111100001111;
20'b00010110000110011011: color_data = 12'b111100001111;
20'b00010110000110011100: color_data = 12'b111100001111;
20'b00010110000110011101: color_data = 12'b111100001111;
20'b00010110000110011110: color_data = 12'b111100001111;
20'b00010110000110011111: color_data = 12'b111100001111;
20'b00010110000110100000: color_data = 12'b111100001111;
20'b00010110000110100001: color_data = 12'b111100001111;
20'b00010110000110100010: color_data = 12'b111100001111;
20'b00010110000110100011: color_data = 12'b111100001111;
20'b00010110000110100100: color_data = 12'b111100001111;
20'b00010110000110100101: color_data = 12'b111100001111;
20'b00010110000110100110: color_data = 12'b111100001111;
20'b00010110000110100111: color_data = 12'b111100001111;
20'b00010110000110101000: color_data = 12'b111100001111;
20'b00010110000110101001: color_data = 12'b111100001111;
20'b00010110000110101010: color_data = 12'b111100001111;
20'b00010110000110101011: color_data = 12'b111100001111;
20'b00010110000110101100: color_data = 12'b111100001111;
20'b00010110000110101101: color_data = 12'b111100001111;
20'b00010110000110101110: color_data = 12'b111100001111;
20'b00010110000110101111: color_data = 12'b111100001111;
20'b00010110000110110000: color_data = 12'b111100001111;
20'b00010110000110110001: color_data = 12'b111100001111;
20'b00010110000110110010: color_data = 12'b111100001111;
20'b00010110000110110011: color_data = 12'b111100001111;
20'b00010110000110110100: color_data = 12'b111100001111;
20'b00010110000110110101: color_data = 12'b111100001111;
20'b00010110000110110110: color_data = 12'b111100001111;
20'b00010110000110110111: color_data = 12'b111100001111;
20'b00010110010011010011: color_data = 12'b000000001111;
20'b00010110010011010100: color_data = 12'b000000001111;
20'b00010110010011010101: color_data = 12'b000000001111;
20'b00010110010011010110: color_data = 12'b000000001111;
20'b00010110010011010111: color_data = 12'b000000001111;
20'b00010110010011011000: color_data = 12'b000000001111;
20'b00010110010011011001: color_data = 12'b000000001111;
20'b00010110010011011010: color_data = 12'b000000001111;
20'b00010110010011011011: color_data = 12'b000000001111;
20'b00010110010011011100: color_data = 12'b000000001111;
20'b00010110010011011101: color_data = 12'b000000001111;
20'b00010110010011011110: color_data = 12'b000000001111;
20'b00010110010011011111: color_data = 12'b000000001111;
20'b00010110010011100000: color_data = 12'b000000001111;
20'b00010110010011100001: color_data = 12'b000000001111;
20'b00010110010011100010: color_data = 12'b000000001111;
20'b00010110010011100011: color_data = 12'b000000001111;
20'b00010110010011100100: color_data = 12'b000000001111;
20'b00010110010011100101: color_data = 12'b000000001111;
20'b00010110010011100110: color_data = 12'b000000001111;
20'b00010110010011100111: color_data = 12'b000000001111;
20'b00010110010011101000: color_data = 12'b000000001111;
20'b00010110010011101001: color_data = 12'b000000001111;
20'b00010110010011101010: color_data = 12'b000000001111;
20'b00010110010011101011: color_data = 12'b000000001111;
20'b00010110010011101100: color_data = 12'b000000001111;
20'b00010110010011101101: color_data = 12'b000000001111;
20'b00010110010011101110: color_data = 12'b000000001111;
20'b00010110010011101111: color_data = 12'b000000001111;
20'b00010110010011110000: color_data = 12'b000000001111;
20'b00010110010011110001: color_data = 12'b000000001111;
20'b00010110010011110010: color_data = 12'b000000001111;
20'b00010110010011110011: color_data = 12'b000000001111;
20'b00010110010011110100: color_data = 12'b000000001111;
20'b00010110010011110101: color_data = 12'b000000001111;
20'b00010110010011110110: color_data = 12'b000000001111;
20'b00010110010011110111: color_data = 12'b000000001111;
20'b00010110010011111000: color_data = 12'b000000001111;
20'b00010110010011111001: color_data = 12'b000000001111;
20'b00010110010011111010: color_data = 12'b000000001111;
20'b00010110010011111011: color_data = 12'b000000001111;
20'b00010110010100000101: color_data = 12'b000001101111;
20'b00010110010100000110: color_data = 12'b000001101111;
20'b00010110010100000111: color_data = 12'b000001101111;
20'b00010110010100001000: color_data = 12'b000001101111;
20'b00010110010100001001: color_data = 12'b000001101111;
20'b00010110010100001010: color_data = 12'b000001101111;
20'b00010110010100001011: color_data = 12'b000001101111;
20'b00010110010100001100: color_data = 12'b000001101111;
20'b00010110010100001101: color_data = 12'b000001101111;
20'b00010110010100001110: color_data = 12'b000001101111;
20'b00010110010100001111: color_data = 12'b000001101111;
20'b00010110010100010000: color_data = 12'b000001101111;
20'b00010110010100010001: color_data = 12'b000001101111;
20'b00010110010100010010: color_data = 12'b000001101111;
20'b00010110010100010011: color_data = 12'b000001101111;
20'b00010110010100010100: color_data = 12'b000001101111;
20'b00010110010100010101: color_data = 12'b000001101111;
20'b00010110010100010110: color_data = 12'b000001101111;
20'b00010110010100010111: color_data = 12'b000001101111;
20'b00010110010100011000: color_data = 12'b000001101111;
20'b00010110010100011001: color_data = 12'b000001101111;
20'b00010110010100011010: color_data = 12'b000001101111;
20'b00010110010100011011: color_data = 12'b000001101111;
20'b00010110010100011100: color_data = 12'b000001101111;
20'b00010110010100011101: color_data = 12'b000001101111;
20'b00010110010100011110: color_data = 12'b000001101111;
20'b00010110010100011111: color_data = 12'b000001101111;
20'b00010110010100100000: color_data = 12'b000001101111;
20'b00010110010100100001: color_data = 12'b000001101111;
20'b00010110010100100010: color_data = 12'b000001101111;
20'b00010110010100100011: color_data = 12'b000001101111;
20'b00010110010100100100: color_data = 12'b000001101111;
20'b00010110010100101101: color_data = 12'b000011111111;
20'b00010110010100101110: color_data = 12'b000011111111;
20'b00010110010100101111: color_data = 12'b000011111111;
20'b00010110010100110000: color_data = 12'b000011111111;
20'b00010110010100110001: color_data = 12'b000011111111;
20'b00010110010100110010: color_data = 12'b000011111111;
20'b00010110010100110011: color_data = 12'b000011111111;
20'b00010110010100110100: color_data = 12'b000011111111;
20'b00010110010100110101: color_data = 12'b000011111111;
20'b00010110010100110110: color_data = 12'b000011111111;
20'b00010110010100110111: color_data = 12'b000011111111;
20'b00010110010100111000: color_data = 12'b000011111111;
20'b00010110010100111001: color_data = 12'b000011111111;
20'b00010110010100111010: color_data = 12'b000011111111;
20'b00010110010100111011: color_data = 12'b000011111111;
20'b00010110010100111100: color_data = 12'b000011111111;
20'b00010110010100111101: color_data = 12'b000011111111;
20'b00010110010100111110: color_data = 12'b000011111111;
20'b00010110010100111111: color_data = 12'b000011111111;
20'b00010110010101000000: color_data = 12'b000011111111;
20'b00010110010101000001: color_data = 12'b000011111111;
20'b00010110010101000010: color_data = 12'b000011111111;
20'b00010110010101000011: color_data = 12'b000011111111;
20'b00010110010101000100: color_data = 12'b000011111111;
20'b00010110010101000101: color_data = 12'b000011111111;
20'b00010110010101000110: color_data = 12'b000011111111;
20'b00010110010101000111: color_data = 12'b000011111111;
20'b00010110010101001000: color_data = 12'b000011111111;
20'b00010110010101001001: color_data = 12'b000011111111;
20'b00010110010101001010: color_data = 12'b000011111111;
20'b00010110010101001011: color_data = 12'b000011111111;
20'b00010110010101001100: color_data = 12'b000011111111;
20'b00010110010101001101: color_data = 12'b000011111111;
20'b00010110010101001110: color_data = 12'b000011111111;
20'b00010110010101001111: color_data = 12'b000011111111;
20'b00010110010101010000: color_data = 12'b000011111111;
20'b00010110010101010001: color_data = 12'b000011111111;
20'b00010110010101010010: color_data = 12'b000011111111;
20'b00010110010101010011: color_data = 12'b000011111111;
20'b00010110010101010100: color_data = 12'b000011111111;
20'b00010110010101010101: color_data = 12'b000011111111;
20'b00010110010101011111: color_data = 12'b111101110000;
20'b00010110010101100000: color_data = 12'b111101110000;
20'b00010110010101100001: color_data = 12'b111101110000;
20'b00010110010101100010: color_data = 12'b111101110000;
20'b00010110010101100011: color_data = 12'b111101110000;
20'b00010110010101100100: color_data = 12'b111101110000;
20'b00010110010101100101: color_data = 12'b111101110000;
20'b00010110010101100110: color_data = 12'b111101110000;
20'b00010110010101100111: color_data = 12'b111101110000;
20'b00010110010101101000: color_data = 12'b111101110000;
20'b00010110010101101001: color_data = 12'b111101110000;
20'b00010110010101101010: color_data = 12'b111101110000;
20'b00010110010101101011: color_data = 12'b111101110000;
20'b00010110010101101100: color_data = 12'b111101110000;
20'b00010110010101101101: color_data = 12'b111101110000;
20'b00010110010101101110: color_data = 12'b111101110000;
20'b00010110010101101111: color_data = 12'b111101110000;
20'b00010110010101110000: color_data = 12'b111101110000;
20'b00010110010101110001: color_data = 12'b111101110000;
20'b00010110010101110010: color_data = 12'b111101110000;
20'b00010110010101110011: color_data = 12'b111101110000;
20'b00010110010101110100: color_data = 12'b111101110000;
20'b00010110010101110101: color_data = 12'b111101110000;
20'b00010110010101110110: color_data = 12'b111101110000;
20'b00010110010101110111: color_data = 12'b111101110000;
20'b00010110010101111000: color_data = 12'b111101110000;
20'b00010110010101111001: color_data = 12'b111101110000;
20'b00010110010101111010: color_data = 12'b111101110000;
20'b00010110010101111011: color_data = 12'b111101110000;
20'b00010110010101111100: color_data = 12'b111101110000;
20'b00010110010101111101: color_data = 12'b111101110000;
20'b00010110010101111110: color_data = 12'b111101110000;
20'b00010110010110000111: color_data = 12'b000011110000;
20'b00010110010110001000: color_data = 12'b000011110000;
20'b00010110010110001001: color_data = 12'b000011110000;
20'b00010110010110001010: color_data = 12'b000011110000;
20'b00010110010110001011: color_data = 12'b000011110000;
20'b00010110010110001100: color_data = 12'b000011110000;
20'b00010110010110001101: color_data = 12'b000011110000;
20'b00010110010110001110: color_data = 12'b000011110000;
20'b00010110010110001111: color_data = 12'b000011110000;
20'b00010110010110011000: color_data = 12'b111100001111;
20'b00010110010110011001: color_data = 12'b111100001111;
20'b00010110010110011010: color_data = 12'b111100001111;
20'b00010110010110011011: color_data = 12'b111100001111;
20'b00010110010110011100: color_data = 12'b111100001111;
20'b00010110010110011101: color_data = 12'b111100001111;
20'b00010110010110011110: color_data = 12'b111100001111;
20'b00010110010110011111: color_data = 12'b111100001111;
20'b00010110010110100000: color_data = 12'b111100001111;
20'b00010110010110100001: color_data = 12'b111100001111;
20'b00010110010110100010: color_data = 12'b111100001111;
20'b00010110010110100011: color_data = 12'b111100001111;
20'b00010110010110100100: color_data = 12'b111100001111;
20'b00010110010110100101: color_data = 12'b111100001111;
20'b00010110010110100110: color_data = 12'b111100001111;
20'b00010110010110100111: color_data = 12'b111100001111;
20'b00010110010110101000: color_data = 12'b111100001111;
20'b00010110010110101001: color_data = 12'b111100001111;
20'b00010110010110101010: color_data = 12'b111100001111;
20'b00010110010110101011: color_data = 12'b111100001111;
20'b00010110010110101100: color_data = 12'b111100001111;
20'b00010110010110101101: color_data = 12'b111100001111;
20'b00010110010110101110: color_data = 12'b111100001111;
20'b00010110010110101111: color_data = 12'b111100001111;
20'b00010110010110110000: color_data = 12'b111100001111;
20'b00010110010110110001: color_data = 12'b111100001111;
20'b00010110010110110010: color_data = 12'b111100001111;
20'b00010110010110110011: color_data = 12'b111100001111;
20'b00010110010110110100: color_data = 12'b111100001111;
20'b00010110010110110101: color_data = 12'b111100001111;
20'b00010110010110110110: color_data = 12'b111100001111;
20'b00010110010110110111: color_data = 12'b111100001111;
20'b00010110100011010011: color_data = 12'b000000001111;
20'b00010110100011010100: color_data = 12'b000000001111;
20'b00010110100011010101: color_data = 12'b000000001111;
20'b00010110100011010110: color_data = 12'b000000001111;
20'b00010110100011010111: color_data = 12'b000000001111;
20'b00010110100011011000: color_data = 12'b000000001111;
20'b00010110100011011001: color_data = 12'b000000001111;
20'b00010110100011011010: color_data = 12'b000000001111;
20'b00010110100011011011: color_data = 12'b000000001111;
20'b00010110100011011100: color_data = 12'b000000001111;
20'b00010110100011011101: color_data = 12'b000000001111;
20'b00010110100011011110: color_data = 12'b000000001111;
20'b00010110100011011111: color_data = 12'b000000001111;
20'b00010110100011100000: color_data = 12'b000000001111;
20'b00010110100011100001: color_data = 12'b000000001111;
20'b00010110100011100010: color_data = 12'b000000001111;
20'b00010110100011100011: color_data = 12'b000000001111;
20'b00010110100011100100: color_data = 12'b000000001111;
20'b00010110100011100101: color_data = 12'b000000001111;
20'b00010110100011100110: color_data = 12'b000000001111;
20'b00010110100011100111: color_data = 12'b000000001111;
20'b00010110100011101000: color_data = 12'b000000001111;
20'b00010110100011101001: color_data = 12'b000000001111;
20'b00010110100011101010: color_data = 12'b000000001111;
20'b00010110100011101011: color_data = 12'b000000001111;
20'b00010110100011101100: color_data = 12'b000000001111;
20'b00010110100011101101: color_data = 12'b000000001111;
20'b00010110100011101110: color_data = 12'b000000001111;
20'b00010110100011101111: color_data = 12'b000000001111;
20'b00010110100011110000: color_data = 12'b000000001111;
20'b00010110100011110001: color_data = 12'b000000001111;
20'b00010110100011110010: color_data = 12'b000000001111;
20'b00010110100011110011: color_data = 12'b000000001111;
20'b00010110100011110100: color_data = 12'b000000001111;
20'b00010110100011110101: color_data = 12'b000000001111;
20'b00010110100011110110: color_data = 12'b000000001111;
20'b00010110100011110111: color_data = 12'b000000001111;
20'b00010110100011111000: color_data = 12'b000000001111;
20'b00010110100011111001: color_data = 12'b000000001111;
20'b00010110100011111010: color_data = 12'b000000001111;
20'b00010110100011111011: color_data = 12'b000000001111;
20'b00010110100100000101: color_data = 12'b000001101111;
20'b00010110100100000110: color_data = 12'b000001101111;
20'b00010110100100000111: color_data = 12'b000001101111;
20'b00010110100100001000: color_data = 12'b000001101111;
20'b00010110100100001001: color_data = 12'b000001101111;
20'b00010110100100001010: color_data = 12'b000001101111;
20'b00010110100100001011: color_data = 12'b000001101111;
20'b00010110100100001100: color_data = 12'b000001101111;
20'b00010110100100001101: color_data = 12'b000001101111;
20'b00010110100100001110: color_data = 12'b000001101111;
20'b00010110100100001111: color_data = 12'b000001101111;
20'b00010110100100010000: color_data = 12'b000001101111;
20'b00010110100100010001: color_data = 12'b000001101111;
20'b00010110100100010010: color_data = 12'b000001101111;
20'b00010110100100010011: color_data = 12'b000001101111;
20'b00010110100100010100: color_data = 12'b000001101111;
20'b00010110100100010101: color_data = 12'b000001101111;
20'b00010110100100010110: color_data = 12'b000001101111;
20'b00010110100100010111: color_data = 12'b000001101111;
20'b00010110100100011000: color_data = 12'b000001101111;
20'b00010110100100011001: color_data = 12'b000001101111;
20'b00010110100100011010: color_data = 12'b000001101111;
20'b00010110100100011011: color_data = 12'b000001101111;
20'b00010110100100011100: color_data = 12'b000001101111;
20'b00010110100100011101: color_data = 12'b000001101111;
20'b00010110100100011110: color_data = 12'b000001101111;
20'b00010110100100011111: color_data = 12'b000001101111;
20'b00010110100100100000: color_data = 12'b000001101111;
20'b00010110100100100001: color_data = 12'b000001101111;
20'b00010110100100100010: color_data = 12'b000001101111;
20'b00010110100100100011: color_data = 12'b000001101111;
20'b00010110100100100100: color_data = 12'b000001101111;
20'b00010110100100101101: color_data = 12'b000011111111;
20'b00010110100100101110: color_data = 12'b000011111111;
20'b00010110100100101111: color_data = 12'b000011111111;
20'b00010110100100110000: color_data = 12'b000011111111;
20'b00010110100100110001: color_data = 12'b000011111111;
20'b00010110100100110010: color_data = 12'b000011111111;
20'b00010110100100110011: color_data = 12'b000011111111;
20'b00010110100100110100: color_data = 12'b000011111111;
20'b00010110100100110101: color_data = 12'b000011111111;
20'b00010110100100110110: color_data = 12'b000011111111;
20'b00010110100100110111: color_data = 12'b000011111111;
20'b00010110100100111000: color_data = 12'b000011111111;
20'b00010110100100111001: color_data = 12'b000011111111;
20'b00010110100100111010: color_data = 12'b000011111111;
20'b00010110100100111011: color_data = 12'b000011111111;
20'b00010110100100111100: color_data = 12'b000011111111;
20'b00010110100100111101: color_data = 12'b000011111111;
20'b00010110100100111110: color_data = 12'b000011111111;
20'b00010110100100111111: color_data = 12'b000011111111;
20'b00010110100101000000: color_data = 12'b000011111111;
20'b00010110100101000001: color_data = 12'b000011111111;
20'b00010110100101000010: color_data = 12'b000011111111;
20'b00010110100101000011: color_data = 12'b000011111111;
20'b00010110100101000100: color_data = 12'b000011111111;
20'b00010110100101000101: color_data = 12'b000011111111;
20'b00010110100101000110: color_data = 12'b000011111111;
20'b00010110100101000111: color_data = 12'b000011111111;
20'b00010110100101001000: color_data = 12'b000011111111;
20'b00010110100101001001: color_data = 12'b000011111111;
20'b00010110100101001010: color_data = 12'b000011111111;
20'b00010110100101001011: color_data = 12'b000011111111;
20'b00010110100101001100: color_data = 12'b000011111111;
20'b00010110100101001101: color_data = 12'b000011111111;
20'b00010110100101001110: color_data = 12'b000011111111;
20'b00010110100101001111: color_data = 12'b000011111111;
20'b00010110100101010000: color_data = 12'b000011111111;
20'b00010110100101010001: color_data = 12'b000011111111;
20'b00010110100101010010: color_data = 12'b000011111111;
20'b00010110100101010011: color_data = 12'b000011111111;
20'b00010110100101010100: color_data = 12'b000011111111;
20'b00010110100101010101: color_data = 12'b000011111111;
20'b00010110100101011111: color_data = 12'b111101110000;
20'b00010110100101100000: color_data = 12'b111101110000;
20'b00010110100101100001: color_data = 12'b111101110000;
20'b00010110100101100010: color_data = 12'b111101110000;
20'b00010110100101100011: color_data = 12'b111101110000;
20'b00010110100101100100: color_data = 12'b111101110000;
20'b00010110100101100101: color_data = 12'b111101110000;
20'b00010110100101100110: color_data = 12'b111101110000;
20'b00010110100101100111: color_data = 12'b111101110000;
20'b00010110100101101000: color_data = 12'b111101110000;
20'b00010110100101101001: color_data = 12'b111101110000;
20'b00010110100101101010: color_data = 12'b111101110000;
20'b00010110100101101011: color_data = 12'b111101110000;
20'b00010110100101101100: color_data = 12'b111101110000;
20'b00010110100101101101: color_data = 12'b111101110000;
20'b00010110100101101110: color_data = 12'b111101110000;
20'b00010110100101101111: color_data = 12'b111101110000;
20'b00010110100101110000: color_data = 12'b111101110000;
20'b00010110100101110001: color_data = 12'b111101110000;
20'b00010110100101110010: color_data = 12'b111101110000;
20'b00010110100101110011: color_data = 12'b111101110000;
20'b00010110100101110100: color_data = 12'b111101110000;
20'b00010110100101110101: color_data = 12'b111101110000;
20'b00010110100101110110: color_data = 12'b111101110000;
20'b00010110100101110111: color_data = 12'b111101110000;
20'b00010110100101111000: color_data = 12'b111101110000;
20'b00010110100101111001: color_data = 12'b111101110000;
20'b00010110100101111010: color_data = 12'b111101110000;
20'b00010110100101111011: color_data = 12'b111101110000;
20'b00010110100101111100: color_data = 12'b111101110000;
20'b00010110100101111101: color_data = 12'b111101110000;
20'b00010110100101111110: color_data = 12'b111101110000;
20'b00010110100110000111: color_data = 12'b000011110000;
20'b00010110100110001000: color_data = 12'b000011110000;
20'b00010110100110001001: color_data = 12'b000011110000;
20'b00010110100110001010: color_data = 12'b000011110000;
20'b00010110100110001011: color_data = 12'b000011110000;
20'b00010110100110001100: color_data = 12'b000011110000;
20'b00010110100110001101: color_data = 12'b000011110000;
20'b00010110100110001110: color_data = 12'b000011110000;
20'b00010110100110001111: color_data = 12'b000011110000;
20'b00010110100110011000: color_data = 12'b111100001111;
20'b00010110100110011001: color_data = 12'b111100001111;
20'b00010110100110011010: color_data = 12'b111100001111;
20'b00010110100110011011: color_data = 12'b111100001111;
20'b00010110100110011100: color_data = 12'b111100001111;
20'b00010110100110011101: color_data = 12'b111100001111;
20'b00010110100110011110: color_data = 12'b111100001111;
20'b00010110100110011111: color_data = 12'b111100001111;
20'b00010110100110100000: color_data = 12'b111100001111;
20'b00010110100110100001: color_data = 12'b111100001111;
20'b00010110100110100010: color_data = 12'b111100001111;
20'b00010110100110100011: color_data = 12'b111100001111;
20'b00010110100110100100: color_data = 12'b111100001111;
20'b00010110100110100101: color_data = 12'b111100001111;
20'b00010110100110100110: color_data = 12'b111100001111;
20'b00010110100110100111: color_data = 12'b111100001111;
20'b00010110100110101000: color_data = 12'b111100001111;
20'b00010110100110101001: color_data = 12'b111100001111;
20'b00010110100110101010: color_data = 12'b111100001111;
20'b00010110100110101011: color_data = 12'b111100001111;
20'b00010110100110101100: color_data = 12'b111100001111;
20'b00010110100110101101: color_data = 12'b111100001111;
20'b00010110100110101110: color_data = 12'b111100001111;
20'b00010110100110101111: color_data = 12'b111100001111;
20'b00010110100110110000: color_data = 12'b111100001111;
20'b00010110100110110001: color_data = 12'b111100001111;
20'b00010110100110110010: color_data = 12'b111100001111;
20'b00010110100110110011: color_data = 12'b111100001111;
20'b00010110100110110100: color_data = 12'b111100001111;
20'b00010110100110110101: color_data = 12'b111100001111;
20'b00010110100110110110: color_data = 12'b111100001111;
20'b00010110100110110111: color_data = 12'b111100001111;
20'b00010110110011010011: color_data = 12'b000000001111;
20'b00010110110011010100: color_data = 12'b000000001111;
20'b00010110110011010101: color_data = 12'b000000001111;
20'b00010110110011010110: color_data = 12'b000000001111;
20'b00010110110011010111: color_data = 12'b000000001111;
20'b00010110110011011000: color_data = 12'b000000001111;
20'b00010110110011011001: color_data = 12'b000000001111;
20'b00010110110011011010: color_data = 12'b000000001111;
20'b00010110110011011011: color_data = 12'b000000001111;
20'b00010110110011011100: color_data = 12'b000000001111;
20'b00010110110011011101: color_data = 12'b000000001111;
20'b00010110110011011110: color_data = 12'b000000001111;
20'b00010110110011011111: color_data = 12'b000000001111;
20'b00010110110011100000: color_data = 12'b000000001111;
20'b00010110110011100001: color_data = 12'b000000001111;
20'b00010110110011100010: color_data = 12'b000000001111;
20'b00010110110011100011: color_data = 12'b000000001111;
20'b00010110110011100100: color_data = 12'b000000001111;
20'b00010110110011100101: color_data = 12'b000000001111;
20'b00010110110011100110: color_data = 12'b000000001111;
20'b00010110110011100111: color_data = 12'b000000001111;
20'b00010110110011101000: color_data = 12'b000000001111;
20'b00010110110011101001: color_data = 12'b000000001111;
20'b00010110110011101010: color_data = 12'b000000001111;
20'b00010110110011101011: color_data = 12'b000000001111;
20'b00010110110011101100: color_data = 12'b000000001111;
20'b00010110110011101101: color_data = 12'b000000001111;
20'b00010110110011101110: color_data = 12'b000000001111;
20'b00010110110011101111: color_data = 12'b000000001111;
20'b00010110110011110000: color_data = 12'b000000001111;
20'b00010110110011110001: color_data = 12'b000000001111;
20'b00010110110011110010: color_data = 12'b000000001111;
20'b00010110110011110011: color_data = 12'b000000001111;
20'b00010110110011110100: color_data = 12'b000000001111;
20'b00010110110011110101: color_data = 12'b000000001111;
20'b00010110110011110110: color_data = 12'b000000001111;
20'b00010110110011110111: color_data = 12'b000000001111;
20'b00010110110011111000: color_data = 12'b000000001111;
20'b00010110110011111001: color_data = 12'b000000001111;
20'b00010110110011111010: color_data = 12'b000000001111;
20'b00010110110011111011: color_data = 12'b000000001111;
20'b00010110110100000101: color_data = 12'b000001101111;
20'b00010110110100000110: color_data = 12'b000001101111;
20'b00010110110100000111: color_data = 12'b000001101111;
20'b00010110110100001000: color_data = 12'b000001101111;
20'b00010110110100001001: color_data = 12'b000001101111;
20'b00010110110100001010: color_data = 12'b000001101111;
20'b00010110110100001011: color_data = 12'b000001101111;
20'b00010110110100001100: color_data = 12'b000001101111;
20'b00010110110100001101: color_data = 12'b000001101111;
20'b00010110110100001110: color_data = 12'b000001101111;
20'b00010110110100001111: color_data = 12'b000001101111;
20'b00010110110100010000: color_data = 12'b000001101111;
20'b00010110110100010001: color_data = 12'b000001101111;
20'b00010110110100010010: color_data = 12'b000001101111;
20'b00010110110100010011: color_data = 12'b000001101111;
20'b00010110110100010100: color_data = 12'b000001101111;
20'b00010110110100010101: color_data = 12'b000001101111;
20'b00010110110100010110: color_data = 12'b000001101111;
20'b00010110110100010111: color_data = 12'b000001101111;
20'b00010110110100011000: color_data = 12'b000001101111;
20'b00010110110100011001: color_data = 12'b000001101111;
20'b00010110110100011010: color_data = 12'b000001101111;
20'b00010110110100011011: color_data = 12'b000001101111;
20'b00010110110100011100: color_data = 12'b000001101111;
20'b00010110110100011101: color_data = 12'b000001101111;
20'b00010110110100011110: color_data = 12'b000001101111;
20'b00010110110100011111: color_data = 12'b000001101111;
20'b00010110110100100000: color_data = 12'b000001101111;
20'b00010110110100100001: color_data = 12'b000001101111;
20'b00010110110100100010: color_data = 12'b000001101111;
20'b00010110110100100011: color_data = 12'b000001101111;
20'b00010110110100100100: color_data = 12'b000001101111;
20'b00010110110100101101: color_data = 12'b000011111111;
20'b00010110110100101110: color_data = 12'b000011111111;
20'b00010110110100101111: color_data = 12'b000011111111;
20'b00010110110100110000: color_data = 12'b000011111111;
20'b00010110110100110001: color_data = 12'b000011111111;
20'b00010110110100110010: color_data = 12'b000011111111;
20'b00010110110100110011: color_data = 12'b000011111111;
20'b00010110110100110100: color_data = 12'b000011111111;
20'b00010110110100110101: color_data = 12'b000011111111;
20'b00010110110100110110: color_data = 12'b000011111111;
20'b00010110110100110111: color_data = 12'b000011111111;
20'b00010110110100111000: color_data = 12'b000011111111;
20'b00010110110100111001: color_data = 12'b000011111111;
20'b00010110110100111010: color_data = 12'b000011111111;
20'b00010110110100111011: color_data = 12'b000011111111;
20'b00010110110100111100: color_data = 12'b000011111111;
20'b00010110110100111101: color_data = 12'b000011111111;
20'b00010110110100111110: color_data = 12'b000011111111;
20'b00010110110100111111: color_data = 12'b000011111111;
20'b00010110110101000000: color_data = 12'b000011111111;
20'b00010110110101000001: color_data = 12'b000011111111;
20'b00010110110101000010: color_data = 12'b000011111111;
20'b00010110110101000011: color_data = 12'b000011111111;
20'b00010110110101000100: color_data = 12'b000011111111;
20'b00010110110101000101: color_data = 12'b000011111111;
20'b00010110110101000110: color_data = 12'b000011111111;
20'b00010110110101000111: color_data = 12'b000011111111;
20'b00010110110101001000: color_data = 12'b000011111111;
20'b00010110110101001001: color_data = 12'b000011111111;
20'b00010110110101001010: color_data = 12'b000011111111;
20'b00010110110101001011: color_data = 12'b000011111111;
20'b00010110110101001100: color_data = 12'b000011111111;
20'b00010110110101001101: color_data = 12'b000011111111;
20'b00010110110101001110: color_data = 12'b000011111111;
20'b00010110110101001111: color_data = 12'b000011111111;
20'b00010110110101010000: color_data = 12'b000011111111;
20'b00010110110101010001: color_data = 12'b000011111111;
20'b00010110110101010010: color_data = 12'b000011111111;
20'b00010110110101010011: color_data = 12'b000011111111;
20'b00010110110101010100: color_data = 12'b000011111111;
20'b00010110110101010101: color_data = 12'b000011111111;
20'b00010110110101011111: color_data = 12'b111101110000;
20'b00010110110101100000: color_data = 12'b111101110000;
20'b00010110110101100001: color_data = 12'b111101110000;
20'b00010110110101100010: color_data = 12'b111101110000;
20'b00010110110101100011: color_data = 12'b111101110000;
20'b00010110110101100100: color_data = 12'b111101110000;
20'b00010110110101100101: color_data = 12'b111101110000;
20'b00010110110101100110: color_data = 12'b111101110000;
20'b00010110110101100111: color_data = 12'b111101110000;
20'b00010110110101101000: color_data = 12'b111101110000;
20'b00010110110101101001: color_data = 12'b111101110000;
20'b00010110110101101010: color_data = 12'b111101110000;
20'b00010110110101101011: color_data = 12'b111101110000;
20'b00010110110101101100: color_data = 12'b111101110000;
20'b00010110110101101101: color_data = 12'b111101110000;
20'b00010110110101101110: color_data = 12'b111101110000;
20'b00010110110101101111: color_data = 12'b111101110000;
20'b00010110110101110000: color_data = 12'b111101110000;
20'b00010110110101110001: color_data = 12'b111101110000;
20'b00010110110101110010: color_data = 12'b111101110000;
20'b00010110110101110011: color_data = 12'b111101110000;
20'b00010110110101110100: color_data = 12'b111101110000;
20'b00010110110101110101: color_data = 12'b111101110000;
20'b00010110110101110110: color_data = 12'b111101110000;
20'b00010110110101110111: color_data = 12'b111101110000;
20'b00010110110101111000: color_data = 12'b111101110000;
20'b00010110110101111001: color_data = 12'b111101110000;
20'b00010110110101111010: color_data = 12'b111101110000;
20'b00010110110101111011: color_data = 12'b111101110000;
20'b00010110110101111100: color_data = 12'b111101110000;
20'b00010110110101111101: color_data = 12'b111101110000;
20'b00010110110101111110: color_data = 12'b111101110000;
20'b00010110110110000111: color_data = 12'b000011110000;
20'b00010110110110001000: color_data = 12'b000011110000;
20'b00010110110110001001: color_data = 12'b000011110000;
20'b00010110110110001010: color_data = 12'b000011110000;
20'b00010110110110001011: color_data = 12'b000011110000;
20'b00010110110110001100: color_data = 12'b000011110000;
20'b00010110110110001101: color_data = 12'b000011110000;
20'b00010110110110001110: color_data = 12'b000011110000;
20'b00010110110110001111: color_data = 12'b000011110000;
20'b00010110110110011000: color_data = 12'b111100001111;
20'b00010110110110011001: color_data = 12'b111100001111;
20'b00010110110110011010: color_data = 12'b111100001111;
20'b00010110110110011011: color_data = 12'b111100001111;
20'b00010110110110011100: color_data = 12'b111100001111;
20'b00010110110110011101: color_data = 12'b111100001111;
20'b00010110110110011110: color_data = 12'b111100001111;
20'b00010110110110011111: color_data = 12'b111100001111;
20'b00010110110110100000: color_data = 12'b111100001111;
20'b00010110110110100001: color_data = 12'b111100001111;
20'b00010110110110100010: color_data = 12'b111100001111;
20'b00010110110110100011: color_data = 12'b111100001111;
20'b00010110110110100100: color_data = 12'b111100001111;
20'b00010110110110100101: color_data = 12'b111100001111;
20'b00010110110110100110: color_data = 12'b111100001111;
20'b00010110110110100111: color_data = 12'b111100001111;
20'b00010110110110101000: color_data = 12'b111100001111;
20'b00010110110110101001: color_data = 12'b111100001111;
20'b00010110110110101010: color_data = 12'b111100001111;
20'b00010110110110101011: color_data = 12'b111100001111;
20'b00010110110110101100: color_data = 12'b111100001111;
20'b00010110110110101101: color_data = 12'b111100001111;
20'b00010110110110101110: color_data = 12'b111100001111;
20'b00010110110110101111: color_data = 12'b111100001111;
20'b00010110110110110000: color_data = 12'b111100001111;
20'b00010110110110110001: color_data = 12'b111100001111;
20'b00010110110110110010: color_data = 12'b111100001111;
20'b00010110110110110011: color_data = 12'b111100001111;
20'b00010110110110110100: color_data = 12'b111100001111;
20'b00010110110110110101: color_data = 12'b111100001111;
20'b00010110110110110110: color_data = 12'b111100001111;
20'b00010110110110110111: color_data = 12'b111100001111;
20'b00010111000011010011: color_data = 12'b000000001111;
20'b00010111000011010100: color_data = 12'b000000001111;
20'b00010111000011010101: color_data = 12'b000000001111;
20'b00010111000011010110: color_data = 12'b000000001111;
20'b00010111000011010111: color_data = 12'b000000001111;
20'b00010111000011011000: color_data = 12'b000000001111;
20'b00010111000011011001: color_data = 12'b000000001111;
20'b00010111000011011010: color_data = 12'b000000001111;
20'b00010111000011011011: color_data = 12'b000000001111;
20'b00010111000011011100: color_data = 12'b000000001111;
20'b00010111000011011101: color_data = 12'b000000001111;
20'b00010111000011011110: color_data = 12'b000000001111;
20'b00010111000011011111: color_data = 12'b000000001111;
20'b00010111000011100000: color_data = 12'b000000001111;
20'b00010111000011100001: color_data = 12'b000000001111;
20'b00010111000011100010: color_data = 12'b000000001111;
20'b00010111000011100011: color_data = 12'b000000001111;
20'b00010111000011100100: color_data = 12'b000000001111;
20'b00010111000011100101: color_data = 12'b000000001111;
20'b00010111000011100110: color_data = 12'b000000001111;
20'b00010111000011100111: color_data = 12'b000000001111;
20'b00010111000011101000: color_data = 12'b000000001111;
20'b00010111000011101001: color_data = 12'b000000001111;
20'b00010111000011101010: color_data = 12'b000000001111;
20'b00010111000011101011: color_data = 12'b000000001111;
20'b00010111000011101100: color_data = 12'b000000001111;
20'b00010111000011101101: color_data = 12'b000000001111;
20'b00010111000011101110: color_data = 12'b000000001111;
20'b00010111000011101111: color_data = 12'b000000001111;
20'b00010111000011110000: color_data = 12'b000000001111;
20'b00010111000011110001: color_data = 12'b000000001111;
20'b00010111000011110010: color_data = 12'b000000001111;
20'b00010111000011110011: color_data = 12'b000000001111;
20'b00010111000011110100: color_data = 12'b000000001111;
20'b00010111000011110101: color_data = 12'b000000001111;
20'b00010111000011110110: color_data = 12'b000000001111;
20'b00010111000011110111: color_data = 12'b000000001111;
20'b00010111000011111000: color_data = 12'b000000001111;
20'b00010111000011111001: color_data = 12'b000000001111;
20'b00010111000011111010: color_data = 12'b000000001111;
20'b00010111000011111011: color_data = 12'b000000001111;
20'b00010111000100000101: color_data = 12'b000001101111;
20'b00010111000100000110: color_data = 12'b000001101111;
20'b00010111000100000111: color_data = 12'b000001101111;
20'b00010111000100001000: color_data = 12'b000001101111;
20'b00010111000100001001: color_data = 12'b000001101111;
20'b00010111000100001010: color_data = 12'b000001101111;
20'b00010111000100001011: color_data = 12'b000001101111;
20'b00010111000100001100: color_data = 12'b000001101111;
20'b00010111000100001101: color_data = 12'b000001101111;
20'b00010111000100001110: color_data = 12'b000001101111;
20'b00010111000100001111: color_data = 12'b000001101111;
20'b00010111000100010000: color_data = 12'b000001101111;
20'b00010111000100010001: color_data = 12'b000001101111;
20'b00010111000100010010: color_data = 12'b000001101111;
20'b00010111000100010011: color_data = 12'b000001101111;
20'b00010111000100010100: color_data = 12'b000001101111;
20'b00010111000100010101: color_data = 12'b000001101111;
20'b00010111000100010110: color_data = 12'b000001101111;
20'b00010111000100010111: color_data = 12'b000001101111;
20'b00010111000100011000: color_data = 12'b000001101111;
20'b00010111000100011001: color_data = 12'b000001101111;
20'b00010111000100011010: color_data = 12'b000001101111;
20'b00010111000100011011: color_data = 12'b000001101111;
20'b00010111000100011100: color_data = 12'b000001101111;
20'b00010111000100011101: color_data = 12'b000001101111;
20'b00010111000100011110: color_data = 12'b000001101111;
20'b00010111000100011111: color_data = 12'b000001101111;
20'b00010111000100100000: color_data = 12'b000001101111;
20'b00010111000100100001: color_data = 12'b000001101111;
20'b00010111000100100010: color_data = 12'b000001101111;
20'b00010111000100100011: color_data = 12'b000001101111;
20'b00010111000100100100: color_data = 12'b000001101111;
20'b00010111000100101101: color_data = 12'b000011111111;
20'b00010111000100101110: color_data = 12'b000011111111;
20'b00010111000100101111: color_data = 12'b000011111111;
20'b00010111000100110000: color_data = 12'b000011111111;
20'b00010111000100110001: color_data = 12'b000011111111;
20'b00010111000100110010: color_data = 12'b000011111111;
20'b00010111000100110011: color_data = 12'b000011111111;
20'b00010111000100110100: color_data = 12'b000011111111;
20'b00010111000100110101: color_data = 12'b000011111111;
20'b00010111000100110110: color_data = 12'b000011111111;
20'b00010111000100110111: color_data = 12'b000011111111;
20'b00010111000100111000: color_data = 12'b000011111111;
20'b00010111000100111001: color_data = 12'b000011111111;
20'b00010111000100111010: color_data = 12'b000011111111;
20'b00010111000100111011: color_data = 12'b000011111111;
20'b00010111000100111100: color_data = 12'b000011111111;
20'b00010111000100111101: color_data = 12'b000011111111;
20'b00010111000100111110: color_data = 12'b000011111111;
20'b00010111000100111111: color_data = 12'b000011111111;
20'b00010111000101000000: color_data = 12'b000011111111;
20'b00010111000101000001: color_data = 12'b000011111111;
20'b00010111000101000010: color_data = 12'b000011111111;
20'b00010111000101000011: color_data = 12'b000011111111;
20'b00010111000101000100: color_data = 12'b000011111111;
20'b00010111000101000101: color_data = 12'b000011111111;
20'b00010111000101000110: color_data = 12'b000011111111;
20'b00010111000101000111: color_data = 12'b000011111111;
20'b00010111000101001000: color_data = 12'b000011111111;
20'b00010111000101001001: color_data = 12'b000011111111;
20'b00010111000101001010: color_data = 12'b000011111111;
20'b00010111000101001011: color_data = 12'b000011111111;
20'b00010111000101001100: color_data = 12'b000011111111;
20'b00010111000101001101: color_data = 12'b000011111111;
20'b00010111000101001110: color_data = 12'b000011111111;
20'b00010111000101001111: color_data = 12'b000011111111;
20'b00010111000101010000: color_data = 12'b000011111111;
20'b00010111000101010001: color_data = 12'b000011111111;
20'b00010111000101010010: color_data = 12'b000011111111;
20'b00010111000101010011: color_data = 12'b000011111111;
20'b00010111000101010100: color_data = 12'b000011111111;
20'b00010111000101010101: color_data = 12'b000011111111;
20'b00010111000101011111: color_data = 12'b111101110000;
20'b00010111000101100000: color_data = 12'b111101110000;
20'b00010111000101100001: color_data = 12'b111101110000;
20'b00010111000101100010: color_data = 12'b111101110000;
20'b00010111000101100011: color_data = 12'b111101110000;
20'b00010111000101100100: color_data = 12'b111101110000;
20'b00010111000101100101: color_data = 12'b111101110000;
20'b00010111000101100110: color_data = 12'b111101110000;
20'b00010111000101100111: color_data = 12'b111101110000;
20'b00010111000101101000: color_data = 12'b111101110000;
20'b00010111000101101001: color_data = 12'b111101110000;
20'b00010111000101101010: color_data = 12'b111101110000;
20'b00010111000101101011: color_data = 12'b111101110000;
20'b00010111000101101100: color_data = 12'b111101110000;
20'b00010111000101101101: color_data = 12'b111101110000;
20'b00010111000101101110: color_data = 12'b111101110000;
20'b00010111000101101111: color_data = 12'b111101110000;
20'b00010111000101110000: color_data = 12'b111101110000;
20'b00010111000101110001: color_data = 12'b111101110000;
20'b00010111000101110010: color_data = 12'b111101110000;
20'b00010111000101110011: color_data = 12'b111101110000;
20'b00010111000101110100: color_data = 12'b111101110000;
20'b00010111000101110101: color_data = 12'b111101110000;
20'b00010111000101110110: color_data = 12'b111101110000;
20'b00010111000101110111: color_data = 12'b111101110000;
20'b00010111000101111000: color_data = 12'b111101110000;
20'b00010111000101111001: color_data = 12'b111101110000;
20'b00010111000101111010: color_data = 12'b111101110000;
20'b00010111000101111011: color_data = 12'b111101110000;
20'b00010111000101111100: color_data = 12'b111101110000;
20'b00010111000101111101: color_data = 12'b111101110000;
20'b00010111000101111110: color_data = 12'b111101110000;
20'b00010111000110000111: color_data = 12'b000011110000;
20'b00010111000110001000: color_data = 12'b000011110000;
20'b00010111000110001001: color_data = 12'b000011110000;
20'b00010111000110001010: color_data = 12'b000011110000;
20'b00010111000110001011: color_data = 12'b000011110000;
20'b00010111000110001100: color_data = 12'b000011110000;
20'b00010111000110001101: color_data = 12'b000011110000;
20'b00010111000110001110: color_data = 12'b000011110000;
20'b00010111000110001111: color_data = 12'b000011110000;
20'b00010111000110011000: color_data = 12'b111100001111;
20'b00010111000110011001: color_data = 12'b111100001111;
20'b00010111000110011010: color_data = 12'b111100001111;
20'b00010111000110011011: color_data = 12'b111100001111;
20'b00010111000110011100: color_data = 12'b111100001111;
20'b00010111000110011101: color_data = 12'b111100001111;
20'b00010111000110011110: color_data = 12'b111100001111;
20'b00010111000110011111: color_data = 12'b111100001111;
20'b00010111000110100000: color_data = 12'b111100001111;
20'b00010111000110100001: color_data = 12'b111100001111;
20'b00010111000110100010: color_data = 12'b111100001111;
20'b00010111000110100011: color_data = 12'b111100001111;
20'b00010111000110100100: color_data = 12'b111100001111;
20'b00010111000110100101: color_data = 12'b111100001111;
20'b00010111000110100110: color_data = 12'b111100001111;
20'b00010111000110100111: color_data = 12'b111100001111;
20'b00010111000110101000: color_data = 12'b111100001111;
20'b00010111000110101001: color_data = 12'b111100001111;
20'b00010111000110101010: color_data = 12'b111100001111;
20'b00010111000110101011: color_data = 12'b111100001111;
20'b00010111000110101100: color_data = 12'b111100001111;
20'b00010111000110101101: color_data = 12'b111100001111;
20'b00010111000110101110: color_data = 12'b111100001111;
20'b00010111000110101111: color_data = 12'b111100001111;
20'b00010111000110110000: color_data = 12'b111100001111;
20'b00010111000110110001: color_data = 12'b111100001111;
20'b00010111000110110010: color_data = 12'b111100001111;
20'b00010111000110110011: color_data = 12'b111100001111;
20'b00010111000110110100: color_data = 12'b111100001111;
20'b00010111000110110101: color_data = 12'b111100001111;
20'b00010111000110110110: color_data = 12'b111100001111;
20'b00010111000110110111: color_data = 12'b111100001111;
20'b00010111010011100100: color_data = 12'b000000001111;
20'b00010111010011100101: color_data = 12'b000000001111;
20'b00010111010011100110: color_data = 12'b000000001111;
20'b00010111010011100111: color_data = 12'b000000001111;
20'b00010111010011101000: color_data = 12'b000000001111;
20'b00010111010011101001: color_data = 12'b000000001111;
20'b00010111010011101010: color_data = 12'b000000001111;
20'b00010111010011101011: color_data = 12'b000000001111;
20'b00010111010100000101: color_data = 12'b000001101111;
20'b00010111010100000110: color_data = 12'b000001101111;
20'b00010111010100000111: color_data = 12'b000001101111;
20'b00010111010100001000: color_data = 12'b000001101111;
20'b00010111010100001001: color_data = 12'b000001101111;
20'b00010111010100001010: color_data = 12'b000001101111;
20'b00010111010100001011: color_data = 12'b000001101111;
20'b00010111010100001100: color_data = 12'b000001101111;
20'b00010111010100111110: color_data = 12'b000011111111;
20'b00010111010100111111: color_data = 12'b000011111111;
20'b00010111010101000000: color_data = 12'b000011111111;
20'b00010111010101000001: color_data = 12'b000011111111;
20'b00010111010101000010: color_data = 12'b000011111111;
20'b00010111010101000011: color_data = 12'b000011111111;
20'b00010111010101000100: color_data = 12'b000011111111;
20'b00010111010101000101: color_data = 12'b000011111111;
20'b00010111010101011111: color_data = 12'b111101110000;
20'b00010111010101100000: color_data = 12'b111101110000;
20'b00010111010101100001: color_data = 12'b111101110000;
20'b00010111010101100010: color_data = 12'b111101110000;
20'b00010111010101100011: color_data = 12'b111101110000;
20'b00010111010101100100: color_data = 12'b111101110000;
20'b00010111010101100101: color_data = 12'b111101110000;
20'b00010111010101100110: color_data = 12'b111101110000;
20'b00010111010101110111: color_data = 12'b111101110000;
20'b00010111010101111000: color_data = 12'b111101110000;
20'b00010111010101111001: color_data = 12'b111101110000;
20'b00010111010101111010: color_data = 12'b111101110000;
20'b00010111010101111011: color_data = 12'b111101110000;
20'b00010111010101111100: color_data = 12'b111101110000;
20'b00010111010101111101: color_data = 12'b111101110000;
20'b00010111010101111110: color_data = 12'b111101110000;
20'b00010111010110000111: color_data = 12'b000011110000;
20'b00010111010110001000: color_data = 12'b000011110000;
20'b00010111010110001001: color_data = 12'b000011110000;
20'b00010111010110001010: color_data = 12'b000011110000;
20'b00010111010110001011: color_data = 12'b000011110000;
20'b00010111010110001100: color_data = 12'b000011110000;
20'b00010111010110001101: color_data = 12'b000011110000;
20'b00010111010110001110: color_data = 12'b000011110000;
20'b00010111010110001111: color_data = 12'b000011110000;
20'b00010111010110011000: color_data = 12'b111100001111;
20'b00010111010110011001: color_data = 12'b111100001111;
20'b00010111010110011010: color_data = 12'b111100001111;
20'b00010111010110011011: color_data = 12'b111100001111;
20'b00010111010110011100: color_data = 12'b111100001111;
20'b00010111010110011101: color_data = 12'b111100001111;
20'b00010111010110011110: color_data = 12'b111100001111;
20'b00010111010110011111: color_data = 12'b111100001111;
20'b00010111100011100100: color_data = 12'b000000001111;
20'b00010111100011100101: color_data = 12'b000000001111;
20'b00010111100011100110: color_data = 12'b000000001111;
20'b00010111100011100111: color_data = 12'b000000001111;
20'b00010111100011101000: color_data = 12'b000000001111;
20'b00010111100011101001: color_data = 12'b000000001111;
20'b00010111100011101010: color_data = 12'b000000001111;
20'b00010111100011101011: color_data = 12'b000000001111;
20'b00010111100100000101: color_data = 12'b000001101111;
20'b00010111100100000110: color_data = 12'b000001101111;
20'b00010111100100000111: color_data = 12'b000001101111;
20'b00010111100100001000: color_data = 12'b000001101111;
20'b00010111100100001001: color_data = 12'b000001101111;
20'b00010111100100001010: color_data = 12'b000001101111;
20'b00010111100100001011: color_data = 12'b000001101111;
20'b00010111100100001100: color_data = 12'b000001101111;
20'b00010111100100111110: color_data = 12'b000011111111;
20'b00010111100100111111: color_data = 12'b000011111111;
20'b00010111100101000000: color_data = 12'b000011111111;
20'b00010111100101000001: color_data = 12'b000011111111;
20'b00010111100101000010: color_data = 12'b000011111111;
20'b00010111100101000011: color_data = 12'b000011111111;
20'b00010111100101000100: color_data = 12'b000011111111;
20'b00010111100101000101: color_data = 12'b000011111111;
20'b00010111100101011111: color_data = 12'b111101110000;
20'b00010111100101100000: color_data = 12'b111101110000;
20'b00010111100101100001: color_data = 12'b111101110000;
20'b00010111100101100010: color_data = 12'b111101110000;
20'b00010111100101100011: color_data = 12'b111101110000;
20'b00010111100101100100: color_data = 12'b111101110000;
20'b00010111100101100101: color_data = 12'b111101110000;
20'b00010111100101100110: color_data = 12'b111101110000;
20'b00010111100101110111: color_data = 12'b111101110000;
20'b00010111100101111000: color_data = 12'b111101110000;
20'b00010111100101111001: color_data = 12'b111101110000;
20'b00010111100101111010: color_data = 12'b111101110000;
20'b00010111100101111011: color_data = 12'b111101110000;
20'b00010111100101111100: color_data = 12'b111101110000;
20'b00010111100101111101: color_data = 12'b111101110000;
20'b00010111100101111110: color_data = 12'b111101110000;
20'b00010111100110000111: color_data = 12'b000011110000;
20'b00010111100110001000: color_data = 12'b000011110000;
20'b00010111100110001001: color_data = 12'b000011110000;
20'b00010111100110001010: color_data = 12'b000011110000;
20'b00010111100110001011: color_data = 12'b000011110000;
20'b00010111100110001100: color_data = 12'b000011110000;
20'b00010111100110001101: color_data = 12'b000011110000;
20'b00010111100110001110: color_data = 12'b000011110000;
20'b00010111100110001111: color_data = 12'b000011110000;
20'b00010111100110011000: color_data = 12'b111100001111;
20'b00010111100110011001: color_data = 12'b111100001111;
20'b00010111100110011010: color_data = 12'b111100001111;
20'b00010111100110011011: color_data = 12'b111100001111;
20'b00010111100110011100: color_data = 12'b111100001111;
20'b00010111100110011101: color_data = 12'b111100001111;
20'b00010111100110011110: color_data = 12'b111100001111;
20'b00010111100110011111: color_data = 12'b111100001111;
20'b00010111110011100100: color_data = 12'b000000001111;
20'b00010111110011100101: color_data = 12'b000000001111;
20'b00010111110011100110: color_data = 12'b000000001111;
20'b00010111110011100111: color_data = 12'b000000001111;
20'b00010111110011101000: color_data = 12'b000000001111;
20'b00010111110011101001: color_data = 12'b000000001111;
20'b00010111110011101010: color_data = 12'b000000001111;
20'b00010111110011101011: color_data = 12'b000000001111;
20'b00010111110100000101: color_data = 12'b000001101111;
20'b00010111110100000110: color_data = 12'b000001101111;
20'b00010111110100000111: color_data = 12'b000001101111;
20'b00010111110100001000: color_data = 12'b000001101111;
20'b00010111110100001001: color_data = 12'b000001101111;
20'b00010111110100001010: color_data = 12'b000001101111;
20'b00010111110100001011: color_data = 12'b000001101111;
20'b00010111110100001100: color_data = 12'b000001101111;
20'b00010111110100111110: color_data = 12'b000011111111;
20'b00010111110100111111: color_data = 12'b000011111111;
20'b00010111110101000000: color_data = 12'b000011111111;
20'b00010111110101000001: color_data = 12'b000011111111;
20'b00010111110101000010: color_data = 12'b000011111111;
20'b00010111110101000011: color_data = 12'b000011111111;
20'b00010111110101000100: color_data = 12'b000011111111;
20'b00010111110101000101: color_data = 12'b000011111111;
20'b00010111110101011111: color_data = 12'b111101110000;
20'b00010111110101100000: color_data = 12'b111101110000;
20'b00010111110101100001: color_data = 12'b111101110000;
20'b00010111110101100010: color_data = 12'b111101110000;
20'b00010111110101100011: color_data = 12'b111101110000;
20'b00010111110101100100: color_data = 12'b111101110000;
20'b00010111110101100101: color_data = 12'b111101110000;
20'b00010111110101100110: color_data = 12'b111101110000;
20'b00010111110101110111: color_data = 12'b111101110000;
20'b00010111110101111000: color_data = 12'b111101110000;
20'b00010111110101111001: color_data = 12'b111101110000;
20'b00010111110101111010: color_data = 12'b111101110000;
20'b00010111110101111011: color_data = 12'b111101110000;
20'b00010111110101111100: color_data = 12'b111101110000;
20'b00010111110101111101: color_data = 12'b111101110000;
20'b00010111110101111110: color_data = 12'b111101110000;
20'b00010111110110000111: color_data = 12'b000011110000;
20'b00010111110110001000: color_data = 12'b000011110000;
20'b00010111110110001001: color_data = 12'b000011110000;
20'b00010111110110001010: color_data = 12'b000011110000;
20'b00010111110110001011: color_data = 12'b000011110000;
20'b00010111110110001100: color_data = 12'b000011110000;
20'b00010111110110001101: color_data = 12'b000011110000;
20'b00010111110110001110: color_data = 12'b000011110000;
20'b00010111110110001111: color_data = 12'b000011110000;
20'b00010111110110011000: color_data = 12'b111100001111;
20'b00010111110110011001: color_data = 12'b111100001111;
20'b00010111110110011010: color_data = 12'b111100001111;
20'b00010111110110011011: color_data = 12'b111100001111;
20'b00010111110110011100: color_data = 12'b111100001111;
20'b00010111110110011101: color_data = 12'b111100001111;
20'b00010111110110011110: color_data = 12'b111100001111;
20'b00010111110110011111: color_data = 12'b111100001111;
20'b00011000000011100100: color_data = 12'b000000001111;
20'b00011000000011100101: color_data = 12'b000000001111;
20'b00011000000011100110: color_data = 12'b000000001111;
20'b00011000000011100111: color_data = 12'b000000001111;
20'b00011000000011101000: color_data = 12'b000000001111;
20'b00011000000011101001: color_data = 12'b000000001111;
20'b00011000000011101010: color_data = 12'b000000001111;
20'b00011000000011101011: color_data = 12'b000000001111;
20'b00011000000100000101: color_data = 12'b000001101111;
20'b00011000000100000110: color_data = 12'b000001101111;
20'b00011000000100000111: color_data = 12'b000001101111;
20'b00011000000100001000: color_data = 12'b000001101111;
20'b00011000000100001001: color_data = 12'b000001101111;
20'b00011000000100001010: color_data = 12'b000001101111;
20'b00011000000100001011: color_data = 12'b000001101111;
20'b00011000000100001100: color_data = 12'b000001101111;
20'b00011000000100111110: color_data = 12'b000011111111;
20'b00011000000100111111: color_data = 12'b000011111111;
20'b00011000000101000000: color_data = 12'b000011111111;
20'b00011000000101000001: color_data = 12'b000011111111;
20'b00011000000101000010: color_data = 12'b000011111111;
20'b00011000000101000011: color_data = 12'b000011111111;
20'b00011000000101000100: color_data = 12'b000011111111;
20'b00011000000101000101: color_data = 12'b000011111111;
20'b00011000000101011111: color_data = 12'b111101110000;
20'b00011000000101100000: color_data = 12'b111101110000;
20'b00011000000101100001: color_data = 12'b111101110000;
20'b00011000000101100010: color_data = 12'b111101110000;
20'b00011000000101100011: color_data = 12'b111101110000;
20'b00011000000101100100: color_data = 12'b111101110000;
20'b00011000000101100101: color_data = 12'b111101110000;
20'b00011000000101100110: color_data = 12'b111101110000;
20'b00011000000101110111: color_data = 12'b111101110000;
20'b00011000000101111000: color_data = 12'b111101110000;
20'b00011000000101111001: color_data = 12'b111101110000;
20'b00011000000101111010: color_data = 12'b111101110000;
20'b00011000000101111011: color_data = 12'b111101110000;
20'b00011000000101111100: color_data = 12'b111101110000;
20'b00011000000101111101: color_data = 12'b111101110000;
20'b00011000000101111110: color_data = 12'b111101110000;
20'b00011000000110000111: color_data = 12'b000011110000;
20'b00011000000110001000: color_data = 12'b000011110000;
20'b00011000000110001001: color_data = 12'b000011110000;
20'b00011000000110001010: color_data = 12'b000011110000;
20'b00011000000110001011: color_data = 12'b000011110000;
20'b00011000000110001100: color_data = 12'b000011110000;
20'b00011000000110001101: color_data = 12'b000011110000;
20'b00011000000110001110: color_data = 12'b000011110000;
20'b00011000000110001111: color_data = 12'b000011110000;
20'b00011000000110011000: color_data = 12'b111100001111;
20'b00011000000110011001: color_data = 12'b111100001111;
20'b00011000000110011010: color_data = 12'b111100001111;
20'b00011000000110011011: color_data = 12'b111100001111;
20'b00011000000110011100: color_data = 12'b111100001111;
20'b00011000000110011101: color_data = 12'b111100001111;
20'b00011000000110011110: color_data = 12'b111100001111;
20'b00011000000110011111: color_data = 12'b111100001111;
20'b00011000010011100100: color_data = 12'b000000001111;
20'b00011000010011100101: color_data = 12'b000000001111;
20'b00011000010011100110: color_data = 12'b000000001111;
20'b00011000010011100111: color_data = 12'b000000001111;
20'b00011000010011101000: color_data = 12'b000000001111;
20'b00011000010011101001: color_data = 12'b000000001111;
20'b00011000010011101010: color_data = 12'b000000001111;
20'b00011000010011101011: color_data = 12'b000000001111;
20'b00011000010100000101: color_data = 12'b000001101111;
20'b00011000010100000110: color_data = 12'b000001101111;
20'b00011000010100000111: color_data = 12'b000001101111;
20'b00011000010100001000: color_data = 12'b000001101111;
20'b00011000010100001001: color_data = 12'b000001101111;
20'b00011000010100001010: color_data = 12'b000001101111;
20'b00011000010100001011: color_data = 12'b000001101111;
20'b00011000010100001100: color_data = 12'b000001101111;
20'b00011000010100111110: color_data = 12'b000011111111;
20'b00011000010100111111: color_data = 12'b000011111111;
20'b00011000010101000000: color_data = 12'b000011111111;
20'b00011000010101000001: color_data = 12'b000011111111;
20'b00011000010101000010: color_data = 12'b000011111111;
20'b00011000010101000011: color_data = 12'b000011111111;
20'b00011000010101000100: color_data = 12'b000011111111;
20'b00011000010101000101: color_data = 12'b000011111111;
20'b00011000010101011111: color_data = 12'b111101110000;
20'b00011000010101100000: color_data = 12'b111101110000;
20'b00011000010101100001: color_data = 12'b111101110000;
20'b00011000010101100010: color_data = 12'b111101110000;
20'b00011000010101100011: color_data = 12'b111101110000;
20'b00011000010101100100: color_data = 12'b111101110000;
20'b00011000010101100101: color_data = 12'b111101110000;
20'b00011000010101100110: color_data = 12'b111101110000;
20'b00011000010101110111: color_data = 12'b111101110000;
20'b00011000010101111000: color_data = 12'b111101110000;
20'b00011000010101111001: color_data = 12'b111101110000;
20'b00011000010101111010: color_data = 12'b111101110000;
20'b00011000010101111011: color_data = 12'b111101110000;
20'b00011000010101111100: color_data = 12'b111101110000;
20'b00011000010101111101: color_data = 12'b111101110000;
20'b00011000010101111110: color_data = 12'b111101110000;
20'b00011000010110000111: color_data = 12'b000011110000;
20'b00011000010110001000: color_data = 12'b000011110000;
20'b00011000010110001001: color_data = 12'b000011110000;
20'b00011000010110001010: color_data = 12'b000011110000;
20'b00011000010110001011: color_data = 12'b000011110000;
20'b00011000010110001100: color_data = 12'b000011110000;
20'b00011000010110001101: color_data = 12'b000011110000;
20'b00011000010110001110: color_data = 12'b000011110000;
20'b00011000010110001111: color_data = 12'b000011110000;
20'b00011000010110011000: color_data = 12'b111100001111;
20'b00011000010110011001: color_data = 12'b111100001111;
20'b00011000010110011010: color_data = 12'b111100001111;
20'b00011000010110011011: color_data = 12'b111100001111;
20'b00011000010110011100: color_data = 12'b111100001111;
20'b00011000010110011101: color_data = 12'b111100001111;
20'b00011000010110011110: color_data = 12'b111100001111;
20'b00011000010110011111: color_data = 12'b111100001111;
20'b00011000100011100100: color_data = 12'b000000001111;
20'b00011000100011100101: color_data = 12'b000000001111;
20'b00011000100011100110: color_data = 12'b000000001111;
20'b00011000100011100111: color_data = 12'b000000001111;
20'b00011000100011101000: color_data = 12'b000000001111;
20'b00011000100011101001: color_data = 12'b000000001111;
20'b00011000100011101010: color_data = 12'b000000001111;
20'b00011000100011101011: color_data = 12'b000000001111;
20'b00011000100100000101: color_data = 12'b000001101111;
20'b00011000100100000110: color_data = 12'b000001101111;
20'b00011000100100000111: color_data = 12'b000001101111;
20'b00011000100100001000: color_data = 12'b000001101111;
20'b00011000100100001001: color_data = 12'b000001101111;
20'b00011000100100001010: color_data = 12'b000001101111;
20'b00011000100100001011: color_data = 12'b000001101111;
20'b00011000100100001100: color_data = 12'b000001101111;
20'b00011000100100111110: color_data = 12'b000011111111;
20'b00011000100100111111: color_data = 12'b000011111111;
20'b00011000100101000000: color_data = 12'b000011111111;
20'b00011000100101000001: color_data = 12'b000011111111;
20'b00011000100101000010: color_data = 12'b000011111111;
20'b00011000100101000011: color_data = 12'b000011111111;
20'b00011000100101000100: color_data = 12'b000011111111;
20'b00011000100101000101: color_data = 12'b000011111111;
20'b00011000100101011111: color_data = 12'b111101110000;
20'b00011000100101100000: color_data = 12'b111101110000;
20'b00011000100101100001: color_data = 12'b111101110000;
20'b00011000100101100010: color_data = 12'b111101110000;
20'b00011000100101100011: color_data = 12'b111101110000;
20'b00011000100101100100: color_data = 12'b111101110000;
20'b00011000100101100101: color_data = 12'b111101110000;
20'b00011000100101100110: color_data = 12'b111101110000;
20'b00011000100101110111: color_data = 12'b111101110000;
20'b00011000100101111000: color_data = 12'b111101110000;
20'b00011000100101111001: color_data = 12'b111101110000;
20'b00011000100101111010: color_data = 12'b111101110000;
20'b00011000100101111011: color_data = 12'b111101110000;
20'b00011000100101111100: color_data = 12'b111101110000;
20'b00011000100101111101: color_data = 12'b111101110000;
20'b00011000100101111110: color_data = 12'b111101110000;
20'b00011000100110000111: color_data = 12'b000011110000;
20'b00011000100110001000: color_data = 12'b000011110000;
20'b00011000100110001001: color_data = 12'b000011110000;
20'b00011000100110001010: color_data = 12'b000011110000;
20'b00011000100110001011: color_data = 12'b000011110000;
20'b00011000100110001100: color_data = 12'b000011110000;
20'b00011000100110001101: color_data = 12'b000011110000;
20'b00011000100110001110: color_data = 12'b000011110000;
20'b00011000100110001111: color_data = 12'b000011110000;
20'b00011000100110011000: color_data = 12'b111100001111;
20'b00011000100110011001: color_data = 12'b111100001111;
20'b00011000100110011010: color_data = 12'b111100001111;
20'b00011000100110011011: color_data = 12'b111100001111;
20'b00011000100110011100: color_data = 12'b111100001111;
20'b00011000100110011101: color_data = 12'b111100001111;
20'b00011000100110011110: color_data = 12'b111100001111;
20'b00011000100110011111: color_data = 12'b111100001111;
20'b00011000110011100100: color_data = 12'b000000001111;
20'b00011000110011100101: color_data = 12'b000000001111;
20'b00011000110011100110: color_data = 12'b000000001111;
20'b00011000110011100111: color_data = 12'b000000001111;
20'b00011000110011101000: color_data = 12'b000000001111;
20'b00011000110011101001: color_data = 12'b000000001111;
20'b00011000110011101010: color_data = 12'b000000001111;
20'b00011000110011101011: color_data = 12'b000000001111;
20'b00011000110100000101: color_data = 12'b000001101111;
20'b00011000110100000110: color_data = 12'b000001101111;
20'b00011000110100000111: color_data = 12'b000001101111;
20'b00011000110100001000: color_data = 12'b000001101111;
20'b00011000110100001001: color_data = 12'b000001101111;
20'b00011000110100001010: color_data = 12'b000001101111;
20'b00011000110100001011: color_data = 12'b000001101111;
20'b00011000110100001100: color_data = 12'b000001101111;
20'b00011000110100111110: color_data = 12'b000011111111;
20'b00011000110100111111: color_data = 12'b000011111111;
20'b00011000110101000000: color_data = 12'b000011111111;
20'b00011000110101000001: color_data = 12'b000011111111;
20'b00011000110101000010: color_data = 12'b000011111111;
20'b00011000110101000011: color_data = 12'b000011111111;
20'b00011000110101000100: color_data = 12'b000011111111;
20'b00011000110101000101: color_data = 12'b000011111111;
20'b00011000110101011111: color_data = 12'b111101110000;
20'b00011000110101100000: color_data = 12'b111101110000;
20'b00011000110101100001: color_data = 12'b111101110000;
20'b00011000110101100010: color_data = 12'b111101110000;
20'b00011000110101100011: color_data = 12'b111101110000;
20'b00011000110101100100: color_data = 12'b111101110000;
20'b00011000110101100101: color_data = 12'b111101110000;
20'b00011000110101100110: color_data = 12'b111101110000;
20'b00011000110101110111: color_data = 12'b111101110000;
20'b00011000110101111000: color_data = 12'b111101110000;
20'b00011000110101111001: color_data = 12'b111101110000;
20'b00011000110101111010: color_data = 12'b111101110000;
20'b00011000110101111011: color_data = 12'b111101110000;
20'b00011000110101111100: color_data = 12'b111101110000;
20'b00011000110101111101: color_data = 12'b111101110000;
20'b00011000110101111110: color_data = 12'b111101110000;
20'b00011000110110000111: color_data = 12'b000011110000;
20'b00011000110110001000: color_data = 12'b000011110000;
20'b00011000110110001001: color_data = 12'b000011110000;
20'b00011000110110001010: color_data = 12'b000011110000;
20'b00011000110110001011: color_data = 12'b000011110000;
20'b00011000110110001100: color_data = 12'b000011110000;
20'b00011000110110001101: color_data = 12'b000011110000;
20'b00011000110110001110: color_data = 12'b000011110000;
20'b00011000110110001111: color_data = 12'b000011110000;
20'b00011000110110011000: color_data = 12'b111100001111;
20'b00011000110110011001: color_data = 12'b111100001111;
20'b00011000110110011010: color_data = 12'b111100001111;
20'b00011000110110011011: color_data = 12'b111100001111;
20'b00011000110110011100: color_data = 12'b111100001111;
20'b00011000110110011101: color_data = 12'b111100001111;
20'b00011000110110011110: color_data = 12'b111100001111;
20'b00011000110110011111: color_data = 12'b111100001111;
20'b00011001000011100100: color_data = 12'b000000001111;
20'b00011001000011100101: color_data = 12'b000000001111;
20'b00011001000011100110: color_data = 12'b000000001111;
20'b00011001000011100111: color_data = 12'b000000001111;
20'b00011001000011101000: color_data = 12'b000000001111;
20'b00011001000011101001: color_data = 12'b000000001111;
20'b00011001000011101010: color_data = 12'b000000001111;
20'b00011001000011101011: color_data = 12'b000000001111;
20'b00011001000100000101: color_data = 12'b000001101111;
20'b00011001000100000110: color_data = 12'b000001101111;
20'b00011001000100000111: color_data = 12'b000001101111;
20'b00011001000100001000: color_data = 12'b000001101111;
20'b00011001000100001001: color_data = 12'b000001101111;
20'b00011001000100001010: color_data = 12'b000001101111;
20'b00011001000100001011: color_data = 12'b000001101111;
20'b00011001000100001100: color_data = 12'b000001101111;
20'b00011001000100111110: color_data = 12'b000011111111;
20'b00011001000100111111: color_data = 12'b000011111111;
20'b00011001000101000000: color_data = 12'b000011111111;
20'b00011001000101000001: color_data = 12'b000011111111;
20'b00011001000101000010: color_data = 12'b000011111111;
20'b00011001000101000011: color_data = 12'b000011111111;
20'b00011001000101000100: color_data = 12'b000011111111;
20'b00011001000101000101: color_data = 12'b000011111111;
20'b00011001000101011111: color_data = 12'b111101110000;
20'b00011001000101100000: color_data = 12'b111101110000;
20'b00011001000101100001: color_data = 12'b111101110000;
20'b00011001000101100010: color_data = 12'b111101110000;
20'b00011001000101100011: color_data = 12'b111101110000;
20'b00011001000101100100: color_data = 12'b111101110000;
20'b00011001000101100101: color_data = 12'b111101110000;
20'b00011001000101100110: color_data = 12'b111101110000;
20'b00011001000101110111: color_data = 12'b111101110000;
20'b00011001000101111000: color_data = 12'b111101110000;
20'b00011001000101111001: color_data = 12'b111101110000;
20'b00011001000101111010: color_data = 12'b111101110000;
20'b00011001000101111011: color_data = 12'b111101110000;
20'b00011001000101111100: color_data = 12'b111101110000;
20'b00011001000101111101: color_data = 12'b111101110000;
20'b00011001000101111110: color_data = 12'b111101110000;
20'b00011001000110000111: color_data = 12'b000011110000;
20'b00011001000110001000: color_data = 12'b000011110000;
20'b00011001000110001001: color_data = 12'b000011110000;
20'b00011001000110001010: color_data = 12'b000011110000;
20'b00011001000110001011: color_data = 12'b000011110000;
20'b00011001000110001100: color_data = 12'b000011110000;
20'b00011001000110001101: color_data = 12'b000011110000;
20'b00011001000110001110: color_data = 12'b000011110000;
20'b00011001000110001111: color_data = 12'b000011110000;
20'b00011001000110011000: color_data = 12'b111100001111;
20'b00011001000110011001: color_data = 12'b111100001111;
20'b00011001000110011010: color_data = 12'b111100001111;
20'b00011001000110011011: color_data = 12'b111100001111;
20'b00011001000110011100: color_data = 12'b111100001111;
20'b00011001000110011101: color_data = 12'b111100001111;
20'b00011001000110011110: color_data = 12'b111100001111;
20'b00011001000110011111: color_data = 12'b111100001111;
20'b00011001010011100100: color_data = 12'b000000001111;
20'b00011001010011100101: color_data = 12'b000000001111;
20'b00011001010011100110: color_data = 12'b000000001111;
20'b00011001010011100111: color_data = 12'b000000001111;
20'b00011001010011101000: color_data = 12'b000000001111;
20'b00011001010011101001: color_data = 12'b000000001111;
20'b00011001010011101010: color_data = 12'b000000001111;
20'b00011001010011101011: color_data = 12'b000000001111;
20'b00011001010100000101: color_data = 12'b000001101111;
20'b00011001010100000110: color_data = 12'b000001101111;
20'b00011001010100000111: color_data = 12'b000001101111;
20'b00011001010100001000: color_data = 12'b000001101111;
20'b00011001010100001001: color_data = 12'b000001101111;
20'b00011001010100001010: color_data = 12'b000001101111;
20'b00011001010100001011: color_data = 12'b000001101111;
20'b00011001010100001100: color_data = 12'b000001101111;
20'b00011001010100111110: color_data = 12'b000011111111;
20'b00011001010100111111: color_data = 12'b000011111111;
20'b00011001010101000000: color_data = 12'b000011111111;
20'b00011001010101000001: color_data = 12'b000011111111;
20'b00011001010101000010: color_data = 12'b000011111111;
20'b00011001010101000011: color_data = 12'b000011111111;
20'b00011001010101000100: color_data = 12'b000011111111;
20'b00011001010101000101: color_data = 12'b000011111111;
20'b00011001010101011111: color_data = 12'b111101110000;
20'b00011001010101100000: color_data = 12'b111101110000;
20'b00011001010101100001: color_data = 12'b111101110000;
20'b00011001010101100010: color_data = 12'b111101110000;
20'b00011001010101100011: color_data = 12'b111101110000;
20'b00011001010101100100: color_data = 12'b111101110000;
20'b00011001010101100101: color_data = 12'b111101110000;
20'b00011001010101100110: color_data = 12'b111101110000;
20'b00011001010101110111: color_data = 12'b111101110000;
20'b00011001010101111000: color_data = 12'b111101110000;
20'b00011001010101111001: color_data = 12'b111101110000;
20'b00011001010101111010: color_data = 12'b111101110000;
20'b00011001010101111011: color_data = 12'b111101110000;
20'b00011001010101111100: color_data = 12'b111101110000;
20'b00011001010101111101: color_data = 12'b111101110000;
20'b00011001010101111110: color_data = 12'b111101110000;
20'b00011001010110000111: color_data = 12'b000011110000;
20'b00011001010110001000: color_data = 12'b000011110000;
20'b00011001010110001001: color_data = 12'b000011110000;
20'b00011001010110001010: color_data = 12'b000011110000;
20'b00011001010110001011: color_data = 12'b000011110000;
20'b00011001010110001100: color_data = 12'b000011110000;
20'b00011001010110001101: color_data = 12'b000011110000;
20'b00011001010110001110: color_data = 12'b000011110000;
20'b00011001010110001111: color_data = 12'b000011110000;
20'b00011001010110011000: color_data = 12'b111100001111;
20'b00011001010110011001: color_data = 12'b111100001111;
20'b00011001010110011010: color_data = 12'b111100001111;
20'b00011001010110011011: color_data = 12'b111100001111;
20'b00011001010110011100: color_data = 12'b111100001111;
20'b00011001010110011101: color_data = 12'b111100001111;
20'b00011001010110011110: color_data = 12'b111100001111;
20'b00011001010110011111: color_data = 12'b111100001111;
20'b00011001100011100100: color_data = 12'b000000001111;
20'b00011001100011100101: color_data = 12'b000000001111;
20'b00011001100011100110: color_data = 12'b000000001111;
20'b00011001100011100111: color_data = 12'b000000001111;
20'b00011001100011101000: color_data = 12'b000000001111;
20'b00011001100011101001: color_data = 12'b000000001111;
20'b00011001100011101010: color_data = 12'b000000001111;
20'b00011001100011101011: color_data = 12'b000000001111;
20'b00011001100100000101: color_data = 12'b000001101111;
20'b00011001100100000110: color_data = 12'b000001101111;
20'b00011001100100000111: color_data = 12'b000001101111;
20'b00011001100100001000: color_data = 12'b000001101111;
20'b00011001100100001001: color_data = 12'b000001101111;
20'b00011001100100001010: color_data = 12'b000001101111;
20'b00011001100100001011: color_data = 12'b000001101111;
20'b00011001100100001100: color_data = 12'b000001101111;
20'b00011001100100111110: color_data = 12'b000011111111;
20'b00011001100100111111: color_data = 12'b000011111111;
20'b00011001100101000000: color_data = 12'b000011111111;
20'b00011001100101000001: color_data = 12'b000011111111;
20'b00011001100101000010: color_data = 12'b000011111111;
20'b00011001100101000011: color_data = 12'b000011111111;
20'b00011001100101000100: color_data = 12'b000011111111;
20'b00011001100101000101: color_data = 12'b000011111111;
20'b00011001100101011111: color_data = 12'b111101110000;
20'b00011001100101100000: color_data = 12'b111101110000;
20'b00011001100101100001: color_data = 12'b111101110000;
20'b00011001100101100010: color_data = 12'b111101110000;
20'b00011001100101100011: color_data = 12'b111101110000;
20'b00011001100101100100: color_data = 12'b111101110000;
20'b00011001100101100101: color_data = 12'b111101110000;
20'b00011001100101100110: color_data = 12'b111101110000;
20'b00011001100101110111: color_data = 12'b111101110000;
20'b00011001100101111000: color_data = 12'b111101110000;
20'b00011001100101111001: color_data = 12'b111101110000;
20'b00011001100101111010: color_data = 12'b111101110000;
20'b00011001100101111011: color_data = 12'b111101110000;
20'b00011001100101111100: color_data = 12'b111101110000;
20'b00011001100101111101: color_data = 12'b111101110000;
20'b00011001100101111110: color_data = 12'b111101110000;
20'b00011001100110000111: color_data = 12'b000011110000;
20'b00011001100110001000: color_data = 12'b000011110000;
20'b00011001100110001001: color_data = 12'b000011110000;
20'b00011001100110001010: color_data = 12'b000011110000;
20'b00011001100110001011: color_data = 12'b000011110000;
20'b00011001100110001100: color_data = 12'b000011110000;
20'b00011001100110001101: color_data = 12'b000011110000;
20'b00011001100110001110: color_data = 12'b000011110000;
20'b00011001100110001111: color_data = 12'b000011110000;
20'b00011001100110011000: color_data = 12'b111100001111;
20'b00011001100110011001: color_data = 12'b111100001111;
20'b00011001100110011010: color_data = 12'b111100001111;
20'b00011001100110011011: color_data = 12'b111100001111;
20'b00011001100110011100: color_data = 12'b111100001111;
20'b00011001100110011101: color_data = 12'b111100001111;
20'b00011001100110011110: color_data = 12'b111100001111;
20'b00011001100110011111: color_data = 12'b111100001111;
20'b00011001110011100100: color_data = 12'b000000001111;
20'b00011001110011100101: color_data = 12'b000000001111;
20'b00011001110011100110: color_data = 12'b000000001111;
20'b00011001110011100111: color_data = 12'b000000001111;
20'b00011001110011101000: color_data = 12'b000000001111;
20'b00011001110011101001: color_data = 12'b000000001111;
20'b00011001110011101010: color_data = 12'b000000001111;
20'b00011001110011101011: color_data = 12'b000000001111;
20'b00011001110100000101: color_data = 12'b000001101111;
20'b00011001110100000110: color_data = 12'b000001101111;
20'b00011001110100000111: color_data = 12'b000001101111;
20'b00011001110100001000: color_data = 12'b000001101111;
20'b00011001110100001001: color_data = 12'b000001101111;
20'b00011001110100001010: color_data = 12'b000001101111;
20'b00011001110100001011: color_data = 12'b000001101111;
20'b00011001110100001100: color_data = 12'b000001101111;
20'b00011001110100111110: color_data = 12'b000011111111;
20'b00011001110100111111: color_data = 12'b000011111111;
20'b00011001110101000000: color_data = 12'b000011111111;
20'b00011001110101000001: color_data = 12'b000011111111;
20'b00011001110101000010: color_data = 12'b000011111111;
20'b00011001110101000011: color_data = 12'b000011111111;
20'b00011001110101000100: color_data = 12'b000011111111;
20'b00011001110101000101: color_data = 12'b000011111111;
20'b00011001110101011111: color_data = 12'b111101110000;
20'b00011001110101100000: color_data = 12'b111101110000;
20'b00011001110101100001: color_data = 12'b111101110000;
20'b00011001110101100010: color_data = 12'b111101110000;
20'b00011001110101100011: color_data = 12'b111101110000;
20'b00011001110101100100: color_data = 12'b111101110000;
20'b00011001110101100101: color_data = 12'b111101110000;
20'b00011001110101100110: color_data = 12'b111101110000;
20'b00011001110101110111: color_data = 12'b111101110000;
20'b00011001110101111000: color_data = 12'b111101110000;
20'b00011001110101111001: color_data = 12'b111101110000;
20'b00011001110101111010: color_data = 12'b111101110000;
20'b00011001110101111011: color_data = 12'b111101110000;
20'b00011001110101111100: color_data = 12'b111101110000;
20'b00011001110101111101: color_data = 12'b111101110000;
20'b00011001110101111110: color_data = 12'b111101110000;
20'b00011001110110000111: color_data = 12'b000011110000;
20'b00011001110110001000: color_data = 12'b000011110000;
20'b00011001110110001001: color_data = 12'b000011110000;
20'b00011001110110001010: color_data = 12'b000011110000;
20'b00011001110110001011: color_data = 12'b000011110000;
20'b00011001110110001100: color_data = 12'b000011110000;
20'b00011001110110001101: color_data = 12'b000011110000;
20'b00011001110110001110: color_data = 12'b000011110000;
20'b00011001110110001111: color_data = 12'b000011110000;
20'b00011001110110011000: color_data = 12'b111100001111;
20'b00011001110110011001: color_data = 12'b111100001111;
20'b00011001110110011010: color_data = 12'b111100001111;
20'b00011001110110011011: color_data = 12'b111100001111;
20'b00011001110110011100: color_data = 12'b111100001111;
20'b00011001110110011101: color_data = 12'b111100001111;
20'b00011001110110011110: color_data = 12'b111100001111;
20'b00011001110110011111: color_data = 12'b111100001111;
20'b00011010000011100100: color_data = 12'b000000001111;
20'b00011010000011100101: color_data = 12'b000000001111;
20'b00011010000011100110: color_data = 12'b000000001111;
20'b00011010000011100111: color_data = 12'b000000001111;
20'b00011010000011101000: color_data = 12'b000000001111;
20'b00011010000011101001: color_data = 12'b000000001111;
20'b00011010000011101010: color_data = 12'b000000001111;
20'b00011010000011101011: color_data = 12'b000000001111;
20'b00011010000100000101: color_data = 12'b000001101111;
20'b00011010000100000110: color_data = 12'b000001101111;
20'b00011010000100000111: color_data = 12'b000001101111;
20'b00011010000100001000: color_data = 12'b000001101111;
20'b00011010000100001001: color_data = 12'b000001101111;
20'b00011010000100001010: color_data = 12'b000001101111;
20'b00011010000100001011: color_data = 12'b000001101111;
20'b00011010000100001100: color_data = 12'b000001101111;
20'b00011010000100111110: color_data = 12'b000011111111;
20'b00011010000100111111: color_data = 12'b000011111111;
20'b00011010000101000000: color_data = 12'b000011111111;
20'b00011010000101000001: color_data = 12'b000011111111;
20'b00011010000101000010: color_data = 12'b000011111111;
20'b00011010000101000011: color_data = 12'b000011111111;
20'b00011010000101000100: color_data = 12'b000011111111;
20'b00011010000101000101: color_data = 12'b000011111111;
20'b00011010000101011111: color_data = 12'b111101110000;
20'b00011010000101100000: color_data = 12'b111101110000;
20'b00011010000101100001: color_data = 12'b111101110000;
20'b00011010000101100010: color_data = 12'b111101110000;
20'b00011010000101100011: color_data = 12'b111101110000;
20'b00011010000101100100: color_data = 12'b111101110000;
20'b00011010000101100101: color_data = 12'b111101110000;
20'b00011010000101100110: color_data = 12'b111101110000;
20'b00011010000101110111: color_data = 12'b111101110000;
20'b00011010000101111000: color_data = 12'b111101110000;
20'b00011010000101111001: color_data = 12'b111101110000;
20'b00011010000101111010: color_data = 12'b111101110000;
20'b00011010000101111011: color_data = 12'b111101110000;
20'b00011010000101111100: color_data = 12'b111101110000;
20'b00011010000101111101: color_data = 12'b111101110000;
20'b00011010000101111110: color_data = 12'b111101110000;
20'b00011010000110000111: color_data = 12'b000011110000;
20'b00011010000110001000: color_data = 12'b000011110000;
20'b00011010000110001001: color_data = 12'b000011110000;
20'b00011010000110001010: color_data = 12'b000011110000;
20'b00011010000110001011: color_data = 12'b000011110000;
20'b00011010000110001100: color_data = 12'b000011110000;
20'b00011010000110001101: color_data = 12'b000011110000;
20'b00011010000110001110: color_data = 12'b000011110000;
20'b00011010000110001111: color_data = 12'b000011110000;
20'b00011010000110011000: color_data = 12'b111100001111;
20'b00011010000110011001: color_data = 12'b111100001111;
20'b00011010000110011010: color_data = 12'b111100001111;
20'b00011010000110011011: color_data = 12'b111100001111;
20'b00011010000110011100: color_data = 12'b111100001111;
20'b00011010000110011101: color_data = 12'b111100001111;
20'b00011010000110011110: color_data = 12'b111100001111;
20'b00011010000110011111: color_data = 12'b111100001111;
20'b00011010010011100100: color_data = 12'b000000001111;
20'b00011010010011100101: color_data = 12'b000000001111;
20'b00011010010011100110: color_data = 12'b000000001111;
20'b00011010010011100111: color_data = 12'b000000001111;
20'b00011010010011101000: color_data = 12'b000000001111;
20'b00011010010011101001: color_data = 12'b000000001111;
20'b00011010010011101010: color_data = 12'b000000001111;
20'b00011010010011101011: color_data = 12'b000000001111;
20'b00011010010100000101: color_data = 12'b000001101111;
20'b00011010010100000110: color_data = 12'b000001101111;
20'b00011010010100000111: color_data = 12'b000001101111;
20'b00011010010100001000: color_data = 12'b000001101111;
20'b00011010010100001001: color_data = 12'b000001101111;
20'b00011010010100001010: color_data = 12'b000001101111;
20'b00011010010100001011: color_data = 12'b000001101111;
20'b00011010010100001100: color_data = 12'b000001101111;
20'b00011010010100001101: color_data = 12'b000001101111;
20'b00011010010100001110: color_data = 12'b000001101111;
20'b00011010010100001111: color_data = 12'b000001101111;
20'b00011010010100010000: color_data = 12'b000001101111;
20'b00011010010100010001: color_data = 12'b000001101111;
20'b00011010010100010010: color_data = 12'b000001101111;
20'b00011010010100010011: color_data = 12'b000001101111;
20'b00011010010100010100: color_data = 12'b000001101111;
20'b00011010010100010101: color_data = 12'b000001101111;
20'b00011010010100010110: color_data = 12'b000001101111;
20'b00011010010100010111: color_data = 12'b000001101111;
20'b00011010010100011000: color_data = 12'b000001101111;
20'b00011010010100011001: color_data = 12'b000001101111;
20'b00011010010100011010: color_data = 12'b000001101111;
20'b00011010010100011011: color_data = 12'b000001101111;
20'b00011010010100011100: color_data = 12'b000001101111;
20'b00011010010100011101: color_data = 12'b000001101111;
20'b00011010010100011110: color_data = 12'b000001101111;
20'b00011010010100011111: color_data = 12'b000001101111;
20'b00011010010100100000: color_data = 12'b000001101111;
20'b00011010010100100001: color_data = 12'b000001101111;
20'b00011010010100100010: color_data = 12'b000001101111;
20'b00011010010100100011: color_data = 12'b000001101111;
20'b00011010010100100100: color_data = 12'b000001101111;
20'b00011010010100111110: color_data = 12'b000011111111;
20'b00011010010100111111: color_data = 12'b000011111111;
20'b00011010010101000000: color_data = 12'b000011111111;
20'b00011010010101000001: color_data = 12'b000011111111;
20'b00011010010101000010: color_data = 12'b000011111111;
20'b00011010010101000011: color_data = 12'b000011111111;
20'b00011010010101000100: color_data = 12'b000011111111;
20'b00011010010101000101: color_data = 12'b000011111111;
20'b00011010010101011111: color_data = 12'b111101110000;
20'b00011010010101100000: color_data = 12'b111101110000;
20'b00011010010101100001: color_data = 12'b111101110000;
20'b00011010010101100010: color_data = 12'b111101110000;
20'b00011010010101100011: color_data = 12'b111101110000;
20'b00011010010101100100: color_data = 12'b111101110000;
20'b00011010010101100101: color_data = 12'b111101110000;
20'b00011010010101100110: color_data = 12'b111101110000;
20'b00011010010101100111: color_data = 12'b111101110000;
20'b00011010010101101000: color_data = 12'b111101110000;
20'b00011010010101101001: color_data = 12'b111101110000;
20'b00011010010101101010: color_data = 12'b111101110000;
20'b00011010010101101011: color_data = 12'b111101110000;
20'b00011010010101101100: color_data = 12'b111101110000;
20'b00011010010101101101: color_data = 12'b111101110000;
20'b00011010010101101110: color_data = 12'b111101110000;
20'b00011010010101101111: color_data = 12'b111101110000;
20'b00011010010101110000: color_data = 12'b111101110000;
20'b00011010010101110001: color_data = 12'b111101110000;
20'b00011010010101110010: color_data = 12'b111101110000;
20'b00011010010101110011: color_data = 12'b111101110000;
20'b00011010010101110100: color_data = 12'b111101110000;
20'b00011010010101110101: color_data = 12'b111101110000;
20'b00011010010101110110: color_data = 12'b111101110000;
20'b00011010010110000111: color_data = 12'b000011110000;
20'b00011010010110001000: color_data = 12'b000011110000;
20'b00011010010110001001: color_data = 12'b000011110000;
20'b00011010010110001010: color_data = 12'b000011110000;
20'b00011010010110001011: color_data = 12'b000011110000;
20'b00011010010110001100: color_data = 12'b000011110000;
20'b00011010010110001101: color_data = 12'b000011110000;
20'b00011010010110001110: color_data = 12'b000011110000;
20'b00011010010110001111: color_data = 12'b000011110000;
20'b00011010010110011000: color_data = 12'b111100001111;
20'b00011010010110011001: color_data = 12'b111100001111;
20'b00011010010110011010: color_data = 12'b111100001111;
20'b00011010010110011011: color_data = 12'b111100001111;
20'b00011010010110011100: color_data = 12'b111100001111;
20'b00011010010110011101: color_data = 12'b111100001111;
20'b00011010010110011110: color_data = 12'b111100001111;
20'b00011010010110011111: color_data = 12'b111100001111;
20'b00011010010110100000: color_data = 12'b111100001111;
20'b00011010010110100001: color_data = 12'b111100001111;
20'b00011010010110100010: color_data = 12'b111100001111;
20'b00011010010110100011: color_data = 12'b111100001111;
20'b00011010010110100100: color_data = 12'b111100001111;
20'b00011010010110100101: color_data = 12'b111100001111;
20'b00011010010110100110: color_data = 12'b111100001111;
20'b00011010010110100111: color_data = 12'b111100001111;
20'b00011010010110101000: color_data = 12'b111100001111;
20'b00011010010110101001: color_data = 12'b111100001111;
20'b00011010010110101010: color_data = 12'b111100001111;
20'b00011010010110101011: color_data = 12'b111100001111;
20'b00011010010110101100: color_data = 12'b111100001111;
20'b00011010010110101101: color_data = 12'b111100001111;
20'b00011010010110101110: color_data = 12'b111100001111;
20'b00011010010110101111: color_data = 12'b111100001111;
20'b00011010010110110000: color_data = 12'b111100001111;
20'b00011010010110110001: color_data = 12'b111100001111;
20'b00011010010110110010: color_data = 12'b111100001111;
20'b00011010010110110011: color_data = 12'b111100001111;
20'b00011010010110110100: color_data = 12'b111100001111;
20'b00011010010110110101: color_data = 12'b111100001111;
20'b00011010010110110110: color_data = 12'b111100001111;
20'b00011010010110110111: color_data = 12'b111100001111;
20'b00011010100011100100: color_data = 12'b000000001111;
20'b00011010100011100101: color_data = 12'b000000001111;
20'b00011010100011100110: color_data = 12'b000000001111;
20'b00011010100011100111: color_data = 12'b000000001111;
20'b00011010100011101000: color_data = 12'b000000001111;
20'b00011010100011101001: color_data = 12'b000000001111;
20'b00011010100011101010: color_data = 12'b000000001111;
20'b00011010100011101011: color_data = 12'b000000001111;
20'b00011010100100000101: color_data = 12'b000001101111;
20'b00011010100100000110: color_data = 12'b000001101111;
20'b00011010100100000111: color_data = 12'b000001101111;
20'b00011010100100001000: color_data = 12'b000001101111;
20'b00011010100100001001: color_data = 12'b000001101111;
20'b00011010100100001010: color_data = 12'b000001101111;
20'b00011010100100001011: color_data = 12'b000001101111;
20'b00011010100100001100: color_data = 12'b000001101111;
20'b00011010100100001101: color_data = 12'b000001101111;
20'b00011010100100001110: color_data = 12'b000001101111;
20'b00011010100100001111: color_data = 12'b000001101111;
20'b00011010100100010000: color_data = 12'b000001101111;
20'b00011010100100010001: color_data = 12'b000001101111;
20'b00011010100100010010: color_data = 12'b000001101111;
20'b00011010100100010011: color_data = 12'b000001101111;
20'b00011010100100010100: color_data = 12'b000001101111;
20'b00011010100100010101: color_data = 12'b000001101111;
20'b00011010100100010110: color_data = 12'b000001101111;
20'b00011010100100010111: color_data = 12'b000001101111;
20'b00011010100100011000: color_data = 12'b000001101111;
20'b00011010100100011001: color_data = 12'b000001101111;
20'b00011010100100011010: color_data = 12'b000001101111;
20'b00011010100100011011: color_data = 12'b000001101111;
20'b00011010100100011100: color_data = 12'b000001101111;
20'b00011010100100011101: color_data = 12'b000001101111;
20'b00011010100100011110: color_data = 12'b000001101111;
20'b00011010100100011111: color_data = 12'b000001101111;
20'b00011010100100100000: color_data = 12'b000001101111;
20'b00011010100100100001: color_data = 12'b000001101111;
20'b00011010100100100010: color_data = 12'b000001101111;
20'b00011010100100100011: color_data = 12'b000001101111;
20'b00011010100100100100: color_data = 12'b000001101111;
20'b00011010100100111110: color_data = 12'b000011111111;
20'b00011010100100111111: color_data = 12'b000011111111;
20'b00011010100101000000: color_data = 12'b000011111111;
20'b00011010100101000001: color_data = 12'b000011111111;
20'b00011010100101000010: color_data = 12'b000011111111;
20'b00011010100101000011: color_data = 12'b000011111111;
20'b00011010100101000100: color_data = 12'b000011111111;
20'b00011010100101000101: color_data = 12'b000011111111;
20'b00011010100101011111: color_data = 12'b111101110000;
20'b00011010100101100000: color_data = 12'b111101110000;
20'b00011010100101100001: color_data = 12'b111101110000;
20'b00011010100101100010: color_data = 12'b111101110000;
20'b00011010100101100011: color_data = 12'b111101110000;
20'b00011010100101100100: color_data = 12'b111101110000;
20'b00011010100101100101: color_data = 12'b111101110000;
20'b00011010100101100110: color_data = 12'b111101110000;
20'b00011010100101100111: color_data = 12'b111101110000;
20'b00011010100101101000: color_data = 12'b111101110000;
20'b00011010100101101001: color_data = 12'b111101110000;
20'b00011010100101101010: color_data = 12'b111101110000;
20'b00011010100101101011: color_data = 12'b111101110000;
20'b00011010100101101100: color_data = 12'b111101110000;
20'b00011010100101101101: color_data = 12'b111101110000;
20'b00011010100101101110: color_data = 12'b111101110000;
20'b00011010100101101111: color_data = 12'b111101110000;
20'b00011010100101110000: color_data = 12'b111101110000;
20'b00011010100101110001: color_data = 12'b111101110000;
20'b00011010100101110010: color_data = 12'b111101110000;
20'b00011010100101110011: color_data = 12'b111101110000;
20'b00011010100101110100: color_data = 12'b111101110000;
20'b00011010100101110101: color_data = 12'b111101110000;
20'b00011010100101110110: color_data = 12'b111101110000;
20'b00011010100110000111: color_data = 12'b000011110000;
20'b00011010100110001000: color_data = 12'b000011110000;
20'b00011010100110001001: color_data = 12'b000011110000;
20'b00011010100110001010: color_data = 12'b000011110000;
20'b00011010100110001011: color_data = 12'b000011110000;
20'b00011010100110001100: color_data = 12'b000011110000;
20'b00011010100110001101: color_data = 12'b000011110000;
20'b00011010100110001110: color_data = 12'b000011110000;
20'b00011010100110001111: color_data = 12'b000011110000;
20'b00011010100110011000: color_data = 12'b111100001111;
20'b00011010100110011001: color_data = 12'b111100001111;
20'b00011010100110011010: color_data = 12'b111100001111;
20'b00011010100110011011: color_data = 12'b111100001111;
20'b00011010100110011100: color_data = 12'b111100001111;
20'b00011010100110011101: color_data = 12'b111100001111;
20'b00011010100110011110: color_data = 12'b111100001111;
20'b00011010100110011111: color_data = 12'b111100001111;
20'b00011010100110100000: color_data = 12'b111100001111;
20'b00011010100110100001: color_data = 12'b111100001111;
20'b00011010100110100010: color_data = 12'b111100001111;
20'b00011010100110100011: color_data = 12'b111100001111;
20'b00011010100110100100: color_data = 12'b111100001111;
20'b00011010100110100101: color_data = 12'b111100001111;
20'b00011010100110100110: color_data = 12'b111100001111;
20'b00011010100110100111: color_data = 12'b111100001111;
20'b00011010100110101000: color_data = 12'b111100001111;
20'b00011010100110101001: color_data = 12'b111100001111;
20'b00011010100110101010: color_data = 12'b111100001111;
20'b00011010100110101011: color_data = 12'b111100001111;
20'b00011010100110101100: color_data = 12'b111100001111;
20'b00011010100110101101: color_data = 12'b111100001111;
20'b00011010100110101110: color_data = 12'b111100001111;
20'b00011010100110101111: color_data = 12'b111100001111;
20'b00011010100110110000: color_data = 12'b111100001111;
20'b00011010100110110001: color_data = 12'b111100001111;
20'b00011010100110110010: color_data = 12'b111100001111;
20'b00011010100110110011: color_data = 12'b111100001111;
20'b00011010100110110100: color_data = 12'b111100001111;
20'b00011010100110110101: color_data = 12'b111100001111;
20'b00011010100110110110: color_data = 12'b111100001111;
20'b00011010100110110111: color_data = 12'b111100001111;
20'b00011010110011100100: color_data = 12'b000000001111;
20'b00011010110011100101: color_data = 12'b000000001111;
20'b00011010110011100110: color_data = 12'b000000001111;
20'b00011010110011100111: color_data = 12'b000000001111;
20'b00011010110011101000: color_data = 12'b000000001111;
20'b00011010110011101001: color_data = 12'b000000001111;
20'b00011010110011101010: color_data = 12'b000000001111;
20'b00011010110011101011: color_data = 12'b000000001111;
20'b00011010110100000101: color_data = 12'b000001101111;
20'b00011010110100000110: color_data = 12'b000001101111;
20'b00011010110100000111: color_data = 12'b000001101111;
20'b00011010110100001000: color_data = 12'b000001101111;
20'b00011010110100001001: color_data = 12'b000001101111;
20'b00011010110100001010: color_data = 12'b000001101111;
20'b00011010110100001011: color_data = 12'b000001101111;
20'b00011010110100001100: color_data = 12'b000001101111;
20'b00011010110100001101: color_data = 12'b000001101111;
20'b00011010110100001110: color_data = 12'b000001101111;
20'b00011010110100001111: color_data = 12'b000001101111;
20'b00011010110100010000: color_data = 12'b000001101111;
20'b00011010110100010001: color_data = 12'b000001101111;
20'b00011010110100010010: color_data = 12'b000001101111;
20'b00011010110100010011: color_data = 12'b000001101111;
20'b00011010110100010100: color_data = 12'b000001101111;
20'b00011010110100010101: color_data = 12'b000001101111;
20'b00011010110100010110: color_data = 12'b000001101111;
20'b00011010110100010111: color_data = 12'b000001101111;
20'b00011010110100011000: color_data = 12'b000001101111;
20'b00011010110100011001: color_data = 12'b000001101111;
20'b00011010110100011010: color_data = 12'b000001101111;
20'b00011010110100011011: color_data = 12'b000001101111;
20'b00011010110100011100: color_data = 12'b000001101111;
20'b00011010110100011101: color_data = 12'b000001101111;
20'b00011010110100011110: color_data = 12'b000001101111;
20'b00011010110100011111: color_data = 12'b000001101111;
20'b00011010110100100000: color_data = 12'b000001101111;
20'b00011010110100100001: color_data = 12'b000001101111;
20'b00011010110100100010: color_data = 12'b000001101111;
20'b00011010110100100011: color_data = 12'b000001101111;
20'b00011010110100100100: color_data = 12'b000001101111;
20'b00011010110100111110: color_data = 12'b000011111111;
20'b00011010110100111111: color_data = 12'b000011111111;
20'b00011010110101000000: color_data = 12'b000011111111;
20'b00011010110101000001: color_data = 12'b000011111111;
20'b00011010110101000010: color_data = 12'b000011111111;
20'b00011010110101000011: color_data = 12'b000011111111;
20'b00011010110101000100: color_data = 12'b000011111111;
20'b00011010110101000101: color_data = 12'b000011111111;
20'b00011010110101011111: color_data = 12'b111101110000;
20'b00011010110101100000: color_data = 12'b111101110000;
20'b00011010110101100001: color_data = 12'b111101110000;
20'b00011010110101100010: color_data = 12'b111101110000;
20'b00011010110101100011: color_data = 12'b111101110000;
20'b00011010110101100100: color_data = 12'b111101110000;
20'b00011010110101100101: color_data = 12'b111101110000;
20'b00011010110101100110: color_data = 12'b111101110000;
20'b00011010110101100111: color_data = 12'b111101110000;
20'b00011010110101101000: color_data = 12'b111101110000;
20'b00011010110101101001: color_data = 12'b111101110000;
20'b00011010110101101010: color_data = 12'b111101110000;
20'b00011010110101101011: color_data = 12'b111101110000;
20'b00011010110101101100: color_data = 12'b111101110000;
20'b00011010110101101101: color_data = 12'b111101110000;
20'b00011010110101101110: color_data = 12'b111101110000;
20'b00011010110101101111: color_data = 12'b111101110000;
20'b00011010110101110000: color_data = 12'b111101110000;
20'b00011010110101110001: color_data = 12'b111101110000;
20'b00011010110101110010: color_data = 12'b111101110000;
20'b00011010110101110011: color_data = 12'b111101110000;
20'b00011010110101110100: color_data = 12'b111101110000;
20'b00011010110101110101: color_data = 12'b111101110000;
20'b00011010110101110110: color_data = 12'b111101110000;
20'b00011010110110000111: color_data = 12'b000011110000;
20'b00011010110110001000: color_data = 12'b000011110000;
20'b00011010110110001001: color_data = 12'b000011110000;
20'b00011010110110001010: color_data = 12'b000011110000;
20'b00011010110110001011: color_data = 12'b000011110000;
20'b00011010110110001100: color_data = 12'b000011110000;
20'b00011010110110001101: color_data = 12'b000011110000;
20'b00011010110110001110: color_data = 12'b000011110000;
20'b00011010110110001111: color_data = 12'b000011110000;
20'b00011010110110011000: color_data = 12'b111100001111;
20'b00011010110110011001: color_data = 12'b111100001111;
20'b00011010110110011010: color_data = 12'b111100001111;
20'b00011010110110011011: color_data = 12'b111100001111;
20'b00011010110110011100: color_data = 12'b111100001111;
20'b00011010110110011101: color_data = 12'b111100001111;
20'b00011010110110011110: color_data = 12'b111100001111;
20'b00011010110110011111: color_data = 12'b111100001111;
20'b00011010110110100000: color_data = 12'b111100001111;
20'b00011010110110100001: color_data = 12'b111100001111;
20'b00011010110110100010: color_data = 12'b111100001111;
20'b00011010110110100011: color_data = 12'b111100001111;
20'b00011010110110100100: color_data = 12'b111100001111;
20'b00011010110110100101: color_data = 12'b111100001111;
20'b00011010110110100110: color_data = 12'b111100001111;
20'b00011010110110100111: color_data = 12'b111100001111;
20'b00011010110110101000: color_data = 12'b111100001111;
20'b00011010110110101001: color_data = 12'b111100001111;
20'b00011010110110101010: color_data = 12'b111100001111;
20'b00011010110110101011: color_data = 12'b111100001111;
20'b00011010110110101100: color_data = 12'b111100001111;
20'b00011010110110101101: color_data = 12'b111100001111;
20'b00011010110110101110: color_data = 12'b111100001111;
20'b00011010110110101111: color_data = 12'b111100001111;
20'b00011010110110110000: color_data = 12'b111100001111;
20'b00011010110110110001: color_data = 12'b111100001111;
20'b00011010110110110010: color_data = 12'b111100001111;
20'b00011010110110110011: color_data = 12'b111100001111;
20'b00011010110110110100: color_data = 12'b111100001111;
20'b00011010110110110101: color_data = 12'b111100001111;
20'b00011010110110110110: color_data = 12'b111100001111;
20'b00011010110110110111: color_data = 12'b111100001111;
20'b00011011000011100100: color_data = 12'b000000001111;
20'b00011011000011100101: color_data = 12'b000000001111;
20'b00011011000011100110: color_data = 12'b000000001111;
20'b00011011000011100111: color_data = 12'b000000001111;
20'b00011011000011101000: color_data = 12'b000000001111;
20'b00011011000011101001: color_data = 12'b000000001111;
20'b00011011000011101010: color_data = 12'b000000001111;
20'b00011011000011101011: color_data = 12'b000000001111;
20'b00011011000100000101: color_data = 12'b000001101111;
20'b00011011000100000110: color_data = 12'b000001101111;
20'b00011011000100000111: color_data = 12'b000001101111;
20'b00011011000100001000: color_data = 12'b000001101111;
20'b00011011000100001001: color_data = 12'b000001101111;
20'b00011011000100001010: color_data = 12'b000001101111;
20'b00011011000100001011: color_data = 12'b000001101111;
20'b00011011000100001100: color_data = 12'b000001101111;
20'b00011011000100001101: color_data = 12'b000001101111;
20'b00011011000100001110: color_data = 12'b000001101111;
20'b00011011000100001111: color_data = 12'b000001101111;
20'b00011011000100010000: color_data = 12'b000001101111;
20'b00011011000100010001: color_data = 12'b000001101111;
20'b00011011000100010010: color_data = 12'b000001101111;
20'b00011011000100010011: color_data = 12'b000001101111;
20'b00011011000100010100: color_data = 12'b000001101111;
20'b00011011000100010101: color_data = 12'b000001101111;
20'b00011011000100010110: color_data = 12'b000001101111;
20'b00011011000100010111: color_data = 12'b000001101111;
20'b00011011000100011000: color_data = 12'b000001101111;
20'b00011011000100011001: color_data = 12'b000001101111;
20'b00011011000100011010: color_data = 12'b000001101111;
20'b00011011000100011011: color_data = 12'b000001101111;
20'b00011011000100011100: color_data = 12'b000001101111;
20'b00011011000100011101: color_data = 12'b000001101111;
20'b00011011000100011110: color_data = 12'b000001101111;
20'b00011011000100011111: color_data = 12'b000001101111;
20'b00011011000100100000: color_data = 12'b000001101111;
20'b00011011000100100001: color_data = 12'b000001101111;
20'b00011011000100100010: color_data = 12'b000001101111;
20'b00011011000100100011: color_data = 12'b000001101111;
20'b00011011000100100100: color_data = 12'b000001101111;
20'b00011011000100111110: color_data = 12'b000011111111;
20'b00011011000100111111: color_data = 12'b000011111111;
20'b00011011000101000000: color_data = 12'b000011111111;
20'b00011011000101000001: color_data = 12'b000011111111;
20'b00011011000101000010: color_data = 12'b000011111111;
20'b00011011000101000011: color_data = 12'b000011111111;
20'b00011011000101000100: color_data = 12'b000011111111;
20'b00011011000101000101: color_data = 12'b000011111111;
20'b00011011000101011111: color_data = 12'b111101110000;
20'b00011011000101100000: color_data = 12'b111101110000;
20'b00011011000101100001: color_data = 12'b111101110000;
20'b00011011000101100010: color_data = 12'b111101110000;
20'b00011011000101100011: color_data = 12'b111101110000;
20'b00011011000101100100: color_data = 12'b111101110000;
20'b00011011000101100101: color_data = 12'b111101110000;
20'b00011011000101100110: color_data = 12'b111101110000;
20'b00011011000101100111: color_data = 12'b111101110000;
20'b00011011000101101000: color_data = 12'b111101110000;
20'b00011011000101101001: color_data = 12'b111101110000;
20'b00011011000101101010: color_data = 12'b111101110000;
20'b00011011000101101011: color_data = 12'b111101110000;
20'b00011011000101101100: color_data = 12'b111101110000;
20'b00011011000101101101: color_data = 12'b111101110000;
20'b00011011000101101110: color_data = 12'b111101110000;
20'b00011011000101101111: color_data = 12'b111101110000;
20'b00011011000101110000: color_data = 12'b111101110000;
20'b00011011000101110001: color_data = 12'b111101110000;
20'b00011011000101110010: color_data = 12'b111101110000;
20'b00011011000101110011: color_data = 12'b111101110000;
20'b00011011000101110100: color_data = 12'b111101110000;
20'b00011011000101110101: color_data = 12'b111101110000;
20'b00011011000101110110: color_data = 12'b111101110000;
20'b00011011000110000111: color_data = 12'b000011110000;
20'b00011011000110001000: color_data = 12'b000011110000;
20'b00011011000110001001: color_data = 12'b000011110000;
20'b00011011000110001010: color_data = 12'b000011110000;
20'b00011011000110001011: color_data = 12'b000011110000;
20'b00011011000110001100: color_data = 12'b000011110000;
20'b00011011000110001101: color_data = 12'b000011110000;
20'b00011011000110001110: color_data = 12'b000011110000;
20'b00011011000110001111: color_data = 12'b000011110000;
20'b00011011000110011000: color_data = 12'b111100001111;
20'b00011011000110011001: color_data = 12'b111100001111;
20'b00011011000110011010: color_data = 12'b111100001111;
20'b00011011000110011011: color_data = 12'b111100001111;
20'b00011011000110011100: color_data = 12'b111100001111;
20'b00011011000110011101: color_data = 12'b111100001111;
20'b00011011000110011110: color_data = 12'b111100001111;
20'b00011011000110011111: color_data = 12'b111100001111;
20'b00011011000110100000: color_data = 12'b111100001111;
20'b00011011000110100001: color_data = 12'b111100001111;
20'b00011011000110100010: color_data = 12'b111100001111;
20'b00011011000110100011: color_data = 12'b111100001111;
20'b00011011000110100100: color_data = 12'b111100001111;
20'b00011011000110100101: color_data = 12'b111100001111;
20'b00011011000110100110: color_data = 12'b111100001111;
20'b00011011000110100111: color_data = 12'b111100001111;
20'b00011011000110101000: color_data = 12'b111100001111;
20'b00011011000110101001: color_data = 12'b111100001111;
20'b00011011000110101010: color_data = 12'b111100001111;
20'b00011011000110101011: color_data = 12'b111100001111;
20'b00011011000110101100: color_data = 12'b111100001111;
20'b00011011000110101101: color_data = 12'b111100001111;
20'b00011011000110101110: color_data = 12'b111100001111;
20'b00011011000110101111: color_data = 12'b111100001111;
20'b00011011000110110000: color_data = 12'b111100001111;
20'b00011011000110110001: color_data = 12'b111100001111;
20'b00011011000110110010: color_data = 12'b111100001111;
20'b00011011000110110011: color_data = 12'b111100001111;
20'b00011011000110110100: color_data = 12'b111100001111;
20'b00011011000110110101: color_data = 12'b111100001111;
20'b00011011000110110110: color_data = 12'b111100001111;
20'b00011011000110110111: color_data = 12'b111100001111;
20'b00011011010011100100: color_data = 12'b000000001111;
20'b00011011010011100101: color_data = 12'b000000001111;
20'b00011011010011100110: color_data = 12'b000000001111;
20'b00011011010011100111: color_data = 12'b000000001111;
20'b00011011010011101000: color_data = 12'b000000001111;
20'b00011011010011101001: color_data = 12'b000000001111;
20'b00011011010011101010: color_data = 12'b000000001111;
20'b00011011010011101011: color_data = 12'b000000001111;
20'b00011011010100000101: color_data = 12'b000001101111;
20'b00011011010100000110: color_data = 12'b000001101111;
20'b00011011010100000111: color_data = 12'b000001101111;
20'b00011011010100001000: color_data = 12'b000001101111;
20'b00011011010100001001: color_data = 12'b000001101111;
20'b00011011010100001010: color_data = 12'b000001101111;
20'b00011011010100001011: color_data = 12'b000001101111;
20'b00011011010100001100: color_data = 12'b000001101111;
20'b00011011010100001101: color_data = 12'b000001101111;
20'b00011011010100001110: color_data = 12'b000001101111;
20'b00011011010100001111: color_data = 12'b000001101111;
20'b00011011010100010000: color_data = 12'b000001101111;
20'b00011011010100010001: color_data = 12'b000001101111;
20'b00011011010100010010: color_data = 12'b000001101111;
20'b00011011010100010011: color_data = 12'b000001101111;
20'b00011011010100010100: color_data = 12'b000001101111;
20'b00011011010100010101: color_data = 12'b000001101111;
20'b00011011010100010110: color_data = 12'b000001101111;
20'b00011011010100010111: color_data = 12'b000001101111;
20'b00011011010100011000: color_data = 12'b000001101111;
20'b00011011010100011001: color_data = 12'b000001101111;
20'b00011011010100011010: color_data = 12'b000001101111;
20'b00011011010100011011: color_data = 12'b000001101111;
20'b00011011010100011100: color_data = 12'b000001101111;
20'b00011011010100011101: color_data = 12'b000001101111;
20'b00011011010100011110: color_data = 12'b000001101111;
20'b00011011010100011111: color_data = 12'b000001101111;
20'b00011011010100100000: color_data = 12'b000001101111;
20'b00011011010100100001: color_data = 12'b000001101111;
20'b00011011010100100010: color_data = 12'b000001101111;
20'b00011011010100100011: color_data = 12'b000001101111;
20'b00011011010100100100: color_data = 12'b000001101111;
20'b00011011010100111110: color_data = 12'b000011111111;
20'b00011011010100111111: color_data = 12'b000011111111;
20'b00011011010101000000: color_data = 12'b000011111111;
20'b00011011010101000001: color_data = 12'b000011111111;
20'b00011011010101000010: color_data = 12'b000011111111;
20'b00011011010101000011: color_data = 12'b000011111111;
20'b00011011010101000100: color_data = 12'b000011111111;
20'b00011011010101000101: color_data = 12'b000011111111;
20'b00011011010101011111: color_data = 12'b111101110000;
20'b00011011010101100000: color_data = 12'b111101110000;
20'b00011011010101100001: color_data = 12'b111101110000;
20'b00011011010101100010: color_data = 12'b111101110000;
20'b00011011010101100011: color_data = 12'b111101110000;
20'b00011011010101100100: color_data = 12'b111101110000;
20'b00011011010101100101: color_data = 12'b111101110000;
20'b00011011010101100110: color_data = 12'b111101110000;
20'b00011011010101100111: color_data = 12'b111101110000;
20'b00011011010101101000: color_data = 12'b111101110000;
20'b00011011010101101001: color_data = 12'b111101110000;
20'b00011011010101101010: color_data = 12'b111101110000;
20'b00011011010101101011: color_data = 12'b111101110000;
20'b00011011010101101100: color_data = 12'b111101110000;
20'b00011011010101101101: color_data = 12'b111101110000;
20'b00011011010101101110: color_data = 12'b111101110000;
20'b00011011010101101111: color_data = 12'b111101110000;
20'b00011011010101110000: color_data = 12'b111101110000;
20'b00011011010101110001: color_data = 12'b111101110000;
20'b00011011010101110010: color_data = 12'b111101110000;
20'b00011011010101110011: color_data = 12'b111101110000;
20'b00011011010101110100: color_data = 12'b111101110000;
20'b00011011010101110101: color_data = 12'b111101110000;
20'b00011011010101110110: color_data = 12'b111101110000;
20'b00011011010110000111: color_data = 12'b000011110000;
20'b00011011010110001000: color_data = 12'b000011110000;
20'b00011011010110001001: color_data = 12'b000011110000;
20'b00011011010110001010: color_data = 12'b000011110000;
20'b00011011010110001011: color_data = 12'b000011110000;
20'b00011011010110001100: color_data = 12'b000011110000;
20'b00011011010110001101: color_data = 12'b000011110000;
20'b00011011010110001110: color_data = 12'b000011110000;
20'b00011011010110001111: color_data = 12'b000011110000;
20'b00011011010110011000: color_data = 12'b111100001111;
20'b00011011010110011001: color_data = 12'b111100001111;
20'b00011011010110011010: color_data = 12'b111100001111;
20'b00011011010110011011: color_data = 12'b111100001111;
20'b00011011010110011100: color_data = 12'b111100001111;
20'b00011011010110011101: color_data = 12'b111100001111;
20'b00011011010110011110: color_data = 12'b111100001111;
20'b00011011010110011111: color_data = 12'b111100001111;
20'b00011011010110100000: color_data = 12'b111100001111;
20'b00011011010110100001: color_data = 12'b111100001111;
20'b00011011010110100010: color_data = 12'b111100001111;
20'b00011011010110100011: color_data = 12'b111100001111;
20'b00011011010110100100: color_data = 12'b111100001111;
20'b00011011010110100101: color_data = 12'b111100001111;
20'b00011011010110100110: color_data = 12'b111100001111;
20'b00011011010110100111: color_data = 12'b111100001111;
20'b00011011010110101000: color_data = 12'b111100001111;
20'b00011011010110101001: color_data = 12'b111100001111;
20'b00011011010110101010: color_data = 12'b111100001111;
20'b00011011010110101011: color_data = 12'b111100001111;
20'b00011011010110101100: color_data = 12'b111100001111;
20'b00011011010110101101: color_data = 12'b111100001111;
20'b00011011010110101110: color_data = 12'b111100001111;
20'b00011011010110101111: color_data = 12'b111100001111;
20'b00011011010110110000: color_data = 12'b111100001111;
20'b00011011010110110001: color_data = 12'b111100001111;
20'b00011011010110110010: color_data = 12'b111100001111;
20'b00011011010110110011: color_data = 12'b111100001111;
20'b00011011010110110100: color_data = 12'b111100001111;
20'b00011011010110110101: color_data = 12'b111100001111;
20'b00011011010110110110: color_data = 12'b111100001111;
20'b00011011010110110111: color_data = 12'b111100001111;
20'b00011011100011100100: color_data = 12'b000000001111;
20'b00011011100011100101: color_data = 12'b000000001111;
20'b00011011100011100110: color_data = 12'b000000001111;
20'b00011011100011100111: color_data = 12'b000000001111;
20'b00011011100011101000: color_data = 12'b000000001111;
20'b00011011100011101001: color_data = 12'b000000001111;
20'b00011011100011101010: color_data = 12'b000000001111;
20'b00011011100011101011: color_data = 12'b000000001111;
20'b00011011100100000101: color_data = 12'b000001101111;
20'b00011011100100000110: color_data = 12'b000001101111;
20'b00011011100100000111: color_data = 12'b000001101111;
20'b00011011100100001000: color_data = 12'b000001101111;
20'b00011011100100001001: color_data = 12'b000001101111;
20'b00011011100100001010: color_data = 12'b000001101111;
20'b00011011100100001011: color_data = 12'b000001101111;
20'b00011011100100001100: color_data = 12'b000001101111;
20'b00011011100100001101: color_data = 12'b000001101111;
20'b00011011100100001110: color_data = 12'b000001101111;
20'b00011011100100001111: color_data = 12'b000001101111;
20'b00011011100100010000: color_data = 12'b000001101111;
20'b00011011100100010001: color_data = 12'b000001101111;
20'b00011011100100010010: color_data = 12'b000001101111;
20'b00011011100100010011: color_data = 12'b000001101111;
20'b00011011100100010100: color_data = 12'b000001101111;
20'b00011011100100010101: color_data = 12'b000001101111;
20'b00011011100100010110: color_data = 12'b000001101111;
20'b00011011100100010111: color_data = 12'b000001101111;
20'b00011011100100011000: color_data = 12'b000001101111;
20'b00011011100100011001: color_data = 12'b000001101111;
20'b00011011100100011010: color_data = 12'b000001101111;
20'b00011011100100011011: color_data = 12'b000001101111;
20'b00011011100100011100: color_data = 12'b000001101111;
20'b00011011100100011101: color_data = 12'b000001101111;
20'b00011011100100011110: color_data = 12'b000001101111;
20'b00011011100100011111: color_data = 12'b000001101111;
20'b00011011100100100000: color_data = 12'b000001101111;
20'b00011011100100100001: color_data = 12'b000001101111;
20'b00011011100100100010: color_data = 12'b000001101111;
20'b00011011100100100011: color_data = 12'b000001101111;
20'b00011011100100100100: color_data = 12'b000001101111;
20'b00011011100100111110: color_data = 12'b000011111111;
20'b00011011100100111111: color_data = 12'b000011111111;
20'b00011011100101000000: color_data = 12'b000011111111;
20'b00011011100101000001: color_data = 12'b000011111111;
20'b00011011100101000010: color_data = 12'b000011111111;
20'b00011011100101000011: color_data = 12'b000011111111;
20'b00011011100101000100: color_data = 12'b000011111111;
20'b00011011100101000101: color_data = 12'b000011111111;
20'b00011011100101011111: color_data = 12'b111101110000;
20'b00011011100101100000: color_data = 12'b111101110000;
20'b00011011100101100001: color_data = 12'b111101110000;
20'b00011011100101100010: color_data = 12'b111101110000;
20'b00011011100101100011: color_data = 12'b111101110000;
20'b00011011100101100100: color_data = 12'b111101110000;
20'b00011011100101100101: color_data = 12'b111101110000;
20'b00011011100101100110: color_data = 12'b111101110000;
20'b00011011100101100111: color_data = 12'b111101110000;
20'b00011011100101101000: color_data = 12'b111101110000;
20'b00011011100101101001: color_data = 12'b111101110000;
20'b00011011100101101010: color_data = 12'b111101110000;
20'b00011011100101101011: color_data = 12'b111101110000;
20'b00011011100101101100: color_data = 12'b111101110000;
20'b00011011100101101101: color_data = 12'b111101110000;
20'b00011011100101101110: color_data = 12'b111101110000;
20'b00011011100101101111: color_data = 12'b111101110000;
20'b00011011100101110000: color_data = 12'b111101110000;
20'b00011011100101110001: color_data = 12'b111101110000;
20'b00011011100101110010: color_data = 12'b111101110000;
20'b00011011100101110011: color_data = 12'b111101110000;
20'b00011011100101110100: color_data = 12'b111101110000;
20'b00011011100101110101: color_data = 12'b111101110000;
20'b00011011100101110110: color_data = 12'b111101110000;
20'b00011011100110000111: color_data = 12'b000011110000;
20'b00011011100110001000: color_data = 12'b000011110000;
20'b00011011100110001001: color_data = 12'b000011110000;
20'b00011011100110001010: color_data = 12'b000011110000;
20'b00011011100110001011: color_data = 12'b000011110000;
20'b00011011100110001100: color_data = 12'b000011110000;
20'b00011011100110001101: color_data = 12'b000011110000;
20'b00011011100110001110: color_data = 12'b000011110000;
20'b00011011100110001111: color_data = 12'b000011110000;
20'b00011011100110011000: color_data = 12'b111100001111;
20'b00011011100110011001: color_data = 12'b111100001111;
20'b00011011100110011010: color_data = 12'b111100001111;
20'b00011011100110011011: color_data = 12'b111100001111;
20'b00011011100110011100: color_data = 12'b111100001111;
20'b00011011100110011101: color_data = 12'b111100001111;
20'b00011011100110011110: color_data = 12'b111100001111;
20'b00011011100110011111: color_data = 12'b111100001111;
20'b00011011100110100000: color_data = 12'b111100001111;
20'b00011011100110100001: color_data = 12'b111100001111;
20'b00011011100110100010: color_data = 12'b111100001111;
20'b00011011100110100011: color_data = 12'b111100001111;
20'b00011011100110100100: color_data = 12'b111100001111;
20'b00011011100110100101: color_data = 12'b111100001111;
20'b00011011100110100110: color_data = 12'b111100001111;
20'b00011011100110100111: color_data = 12'b111100001111;
20'b00011011100110101000: color_data = 12'b111100001111;
20'b00011011100110101001: color_data = 12'b111100001111;
20'b00011011100110101010: color_data = 12'b111100001111;
20'b00011011100110101011: color_data = 12'b111100001111;
20'b00011011100110101100: color_data = 12'b111100001111;
20'b00011011100110101101: color_data = 12'b111100001111;
20'b00011011100110101110: color_data = 12'b111100001111;
20'b00011011100110101111: color_data = 12'b111100001111;
20'b00011011100110110000: color_data = 12'b111100001111;
20'b00011011100110110001: color_data = 12'b111100001111;
20'b00011011100110110010: color_data = 12'b111100001111;
20'b00011011100110110011: color_data = 12'b111100001111;
20'b00011011100110110100: color_data = 12'b111100001111;
20'b00011011100110110101: color_data = 12'b111100001111;
20'b00011011100110110110: color_data = 12'b111100001111;
20'b00011011100110110111: color_data = 12'b111100001111;
20'b00011011110011100100: color_data = 12'b000000001111;
20'b00011011110011100101: color_data = 12'b000000001111;
20'b00011011110011100110: color_data = 12'b000000001111;
20'b00011011110011100111: color_data = 12'b000000001111;
20'b00011011110011101000: color_data = 12'b000000001111;
20'b00011011110011101001: color_data = 12'b000000001111;
20'b00011011110011101010: color_data = 12'b000000001111;
20'b00011011110011101011: color_data = 12'b000000001111;
20'b00011011110100000101: color_data = 12'b000001101111;
20'b00011011110100000110: color_data = 12'b000001101111;
20'b00011011110100000111: color_data = 12'b000001101111;
20'b00011011110100001000: color_data = 12'b000001101111;
20'b00011011110100001001: color_data = 12'b000001101111;
20'b00011011110100001010: color_data = 12'b000001101111;
20'b00011011110100001011: color_data = 12'b000001101111;
20'b00011011110100001100: color_data = 12'b000001101111;
20'b00011011110100001101: color_data = 12'b000001101111;
20'b00011011110100001110: color_data = 12'b000001101111;
20'b00011011110100001111: color_data = 12'b000001101111;
20'b00011011110100010000: color_data = 12'b000001101111;
20'b00011011110100010001: color_data = 12'b000001101111;
20'b00011011110100010010: color_data = 12'b000001101111;
20'b00011011110100010011: color_data = 12'b000001101111;
20'b00011011110100010100: color_data = 12'b000001101111;
20'b00011011110100010101: color_data = 12'b000001101111;
20'b00011011110100010110: color_data = 12'b000001101111;
20'b00011011110100010111: color_data = 12'b000001101111;
20'b00011011110100011000: color_data = 12'b000001101111;
20'b00011011110100011001: color_data = 12'b000001101111;
20'b00011011110100011010: color_data = 12'b000001101111;
20'b00011011110100011011: color_data = 12'b000001101111;
20'b00011011110100011100: color_data = 12'b000001101111;
20'b00011011110100011101: color_data = 12'b000001101111;
20'b00011011110100011110: color_data = 12'b000001101111;
20'b00011011110100011111: color_data = 12'b000001101111;
20'b00011011110100100000: color_data = 12'b000001101111;
20'b00011011110100100001: color_data = 12'b000001101111;
20'b00011011110100100010: color_data = 12'b000001101111;
20'b00011011110100100011: color_data = 12'b000001101111;
20'b00011011110100100100: color_data = 12'b000001101111;
20'b00011011110100111110: color_data = 12'b000011111111;
20'b00011011110100111111: color_data = 12'b000011111111;
20'b00011011110101000000: color_data = 12'b000011111111;
20'b00011011110101000001: color_data = 12'b000011111111;
20'b00011011110101000010: color_data = 12'b000011111111;
20'b00011011110101000011: color_data = 12'b000011111111;
20'b00011011110101000100: color_data = 12'b000011111111;
20'b00011011110101000101: color_data = 12'b000011111111;
20'b00011011110101011111: color_data = 12'b111101110000;
20'b00011011110101100000: color_data = 12'b111101110000;
20'b00011011110101100001: color_data = 12'b111101110000;
20'b00011011110101100010: color_data = 12'b111101110000;
20'b00011011110101100011: color_data = 12'b111101110000;
20'b00011011110101100100: color_data = 12'b111101110000;
20'b00011011110101100101: color_data = 12'b111101110000;
20'b00011011110101100110: color_data = 12'b111101110000;
20'b00011011110101100111: color_data = 12'b111101110000;
20'b00011011110101101000: color_data = 12'b111101110000;
20'b00011011110101101001: color_data = 12'b111101110000;
20'b00011011110101101010: color_data = 12'b111101110000;
20'b00011011110101101011: color_data = 12'b111101110000;
20'b00011011110101101100: color_data = 12'b111101110000;
20'b00011011110101101101: color_data = 12'b111101110000;
20'b00011011110101101110: color_data = 12'b111101110000;
20'b00011011110101101111: color_data = 12'b111101110000;
20'b00011011110101110000: color_data = 12'b111101110000;
20'b00011011110101110001: color_data = 12'b111101110000;
20'b00011011110101110010: color_data = 12'b111101110000;
20'b00011011110101110011: color_data = 12'b111101110000;
20'b00011011110101110100: color_data = 12'b111101110000;
20'b00011011110101110101: color_data = 12'b111101110000;
20'b00011011110101110110: color_data = 12'b111101110000;
20'b00011011110110000111: color_data = 12'b000011110000;
20'b00011011110110001000: color_data = 12'b000011110000;
20'b00011011110110001001: color_data = 12'b000011110000;
20'b00011011110110001010: color_data = 12'b000011110000;
20'b00011011110110001011: color_data = 12'b000011110000;
20'b00011011110110001100: color_data = 12'b000011110000;
20'b00011011110110001101: color_data = 12'b000011110000;
20'b00011011110110001110: color_data = 12'b000011110000;
20'b00011011110110001111: color_data = 12'b000011110000;
20'b00011011110110011000: color_data = 12'b111100001111;
20'b00011011110110011001: color_data = 12'b111100001111;
20'b00011011110110011010: color_data = 12'b111100001111;
20'b00011011110110011011: color_data = 12'b111100001111;
20'b00011011110110011100: color_data = 12'b111100001111;
20'b00011011110110011101: color_data = 12'b111100001111;
20'b00011011110110011110: color_data = 12'b111100001111;
20'b00011011110110011111: color_data = 12'b111100001111;
20'b00011011110110100000: color_data = 12'b111100001111;
20'b00011011110110100001: color_data = 12'b111100001111;
20'b00011011110110100010: color_data = 12'b111100001111;
20'b00011011110110100011: color_data = 12'b111100001111;
20'b00011011110110100100: color_data = 12'b111100001111;
20'b00011011110110100101: color_data = 12'b111100001111;
20'b00011011110110100110: color_data = 12'b111100001111;
20'b00011011110110100111: color_data = 12'b111100001111;
20'b00011011110110101000: color_data = 12'b111100001111;
20'b00011011110110101001: color_data = 12'b111100001111;
20'b00011011110110101010: color_data = 12'b111100001111;
20'b00011011110110101011: color_data = 12'b111100001111;
20'b00011011110110101100: color_data = 12'b111100001111;
20'b00011011110110101101: color_data = 12'b111100001111;
20'b00011011110110101110: color_data = 12'b111100001111;
20'b00011011110110101111: color_data = 12'b111100001111;
20'b00011011110110110000: color_data = 12'b111100001111;
20'b00011011110110110001: color_data = 12'b111100001111;
20'b00011011110110110010: color_data = 12'b111100001111;
20'b00011011110110110011: color_data = 12'b111100001111;
20'b00011011110110110100: color_data = 12'b111100001111;
20'b00011011110110110101: color_data = 12'b111100001111;
20'b00011011110110110110: color_data = 12'b111100001111;
20'b00011011110110110111: color_data = 12'b111100001111;
20'b00011100000011100100: color_data = 12'b000000001111;
20'b00011100000011100101: color_data = 12'b000000001111;
20'b00011100000011100110: color_data = 12'b000000001111;
20'b00011100000011100111: color_data = 12'b000000001111;
20'b00011100000011101000: color_data = 12'b000000001111;
20'b00011100000011101001: color_data = 12'b000000001111;
20'b00011100000011101010: color_data = 12'b000000001111;
20'b00011100000011101011: color_data = 12'b000000001111;
20'b00011100000100000101: color_data = 12'b000001101111;
20'b00011100000100000110: color_data = 12'b000001101111;
20'b00011100000100000111: color_data = 12'b000001101111;
20'b00011100000100001000: color_data = 12'b000001101111;
20'b00011100000100001001: color_data = 12'b000001101111;
20'b00011100000100001010: color_data = 12'b000001101111;
20'b00011100000100001011: color_data = 12'b000001101111;
20'b00011100000100001100: color_data = 12'b000001101111;
20'b00011100000100001101: color_data = 12'b000001101111;
20'b00011100000100001110: color_data = 12'b000001101111;
20'b00011100000100001111: color_data = 12'b000001101111;
20'b00011100000100010000: color_data = 12'b000001101111;
20'b00011100000100010001: color_data = 12'b000001101111;
20'b00011100000100010010: color_data = 12'b000001101111;
20'b00011100000100010011: color_data = 12'b000001101111;
20'b00011100000100010100: color_data = 12'b000001101111;
20'b00011100000100010101: color_data = 12'b000001101111;
20'b00011100000100010110: color_data = 12'b000001101111;
20'b00011100000100010111: color_data = 12'b000001101111;
20'b00011100000100011000: color_data = 12'b000001101111;
20'b00011100000100011001: color_data = 12'b000001101111;
20'b00011100000100011010: color_data = 12'b000001101111;
20'b00011100000100011011: color_data = 12'b000001101111;
20'b00011100000100011100: color_data = 12'b000001101111;
20'b00011100000100011101: color_data = 12'b000001101111;
20'b00011100000100011110: color_data = 12'b000001101111;
20'b00011100000100011111: color_data = 12'b000001101111;
20'b00011100000100100000: color_data = 12'b000001101111;
20'b00011100000100100001: color_data = 12'b000001101111;
20'b00011100000100100010: color_data = 12'b000001101111;
20'b00011100000100100011: color_data = 12'b000001101111;
20'b00011100000100100100: color_data = 12'b000001101111;
20'b00011100000100111110: color_data = 12'b000011111111;
20'b00011100000100111111: color_data = 12'b000011111111;
20'b00011100000101000000: color_data = 12'b000011111111;
20'b00011100000101000001: color_data = 12'b000011111111;
20'b00011100000101000010: color_data = 12'b000011111111;
20'b00011100000101000011: color_data = 12'b000011111111;
20'b00011100000101000100: color_data = 12'b000011111111;
20'b00011100000101000101: color_data = 12'b000011111111;
20'b00011100000101011111: color_data = 12'b111101110000;
20'b00011100000101100000: color_data = 12'b111101110000;
20'b00011100000101100001: color_data = 12'b111101110000;
20'b00011100000101100010: color_data = 12'b111101110000;
20'b00011100000101100011: color_data = 12'b111101110000;
20'b00011100000101100100: color_data = 12'b111101110000;
20'b00011100000101100101: color_data = 12'b111101110000;
20'b00011100000101100110: color_data = 12'b111101110000;
20'b00011100000101100111: color_data = 12'b111101110000;
20'b00011100000101101000: color_data = 12'b111101110000;
20'b00011100000101101001: color_data = 12'b111101110000;
20'b00011100000101101010: color_data = 12'b111101110000;
20'b00011100000101101011: color_data = 12'b111101110000;
20'b00011100000101101100: color_data = 12'b111101110000;
20'b00011100000101101101: color_data = 12'b111101110000;
20'b00011100000101101110: color_data = 12'b111101110000;
20'b00011100000101101111: color_data = 12'b111101110000;
20'b00011100000101110000: color_data = 12'b111101110000;
20'b00011100000101110001: color_data = 12'b111101110000;
20'b00011100000101110010: color_data = 12'b111101110000;
20'b00011100000101110011: color_data = 12'b111101110000;
20'b00011100000101110100: color_data = 12'b111101110000;
20'b00011100000101110101: color_data = 12'b111101110000;
20'b00011100000101110110: color_data = 12'b111101110000;
20'b00011100000110000111: color_data = 12'b000011110000;
20'b00011100000110001000: color_data = 12'b000011110000;
20'b00011100000110001001: color_data = 12'b000011110000;
20'b00011100000110001010: color_data = 12'b000011110000;
20'b00011100000110001011: color_data = 12'b000011110000;
20'b00011100000110001100: color_data = 12'b000011110000;
20'b00011100000110001101: color_data = 12'b000011110000;
20'b00011100000110001110: color_data = 12'b000011110000;
20'b00011100000110001111: color_data = 12'b000011110000;
20'b00011100000110011000: color_data = 12'b111100001111;
20'b00011100000110011001: color_data = 12'b111100001111;
20'b00011100000110011010: color_data = 12'b111100001111;
20'b00011100000110011011: color_data = 12'b111100001111;
20'b00011100000110011100: color_data = 12'b111100001111;
20'b00011100000110011101: color_data = 12'b111100001111;
20'b00011100000110011110: color_data = 12'b111100001111;
20'b00011100000110011111: color_data = 12'b111100001111;
20'b00011100000110100000: color_data = 12'b111100001111;
20'b00011100000110100001: color_data = 12'b111100001111;
20'b00011100000110100010: color_data = 12'b111100001111;
20'b00011100000110100011: color_data = 12'b111100001111;
20'b00011100000110100100: color_data = 12'b111100001111;
20'b00011100000110100101: color_data = 12'b111100001111;
20'b00011100000110100110: color_data = 12'b111100001111;
20'b00011100000110100111: color_data = 12'b111100001111;
20'b00011100000110101000: color_data = 12'b111100001111;
20'b00011100000110101001: color_data = 12'b111100001111;
20'b00011100000110101010: color_data = 12'b111100001111;
20'b00011100000110101011: color_data = 12'b111100001111;
20'b00011100000110101100: color_data = 12'b111100001111;
20'b00011100000110101101: color_data = 12'b111100001111;
20'b00011100000110101110: color_data = 12'b111100001111;
20'b00011100000110101111: color_data = 12'b111100001111;
20'b00011100000110110000: color_data = 12'b111100001111;
20'b00011100000110110001: color_data = 12'b111100001111;
20'b00011100000110110010: color_data = 12'b111100001111;
20'b00011100000110110011: color_data = 12'b111100001111;
20'b00011100000110110100: color_data = 12'b111100001111;
20'b00011100000110110101: color_data = 12'b111100001111;
20'b00011100000110110110: color_data = 12'b111100001111;
20'b00011100000110110111: color_data = 12'b111100001111;
20'b00011100010011100100: color_data = 12'b000000001111;
20'b00011100010011100101: color_data = 12'b000000001111;
20'b00011100010011100110: color_data = 12'b000000001111;
20'b00011100010011100111: color_data = 12'b000000001111;
20'b00011100010011101000: color_data = 12'b000000001111;
20'b00011100010011101001: color_data = 12'b000000001111;
20'b00011100010011101010: color_data = 12'b000000001111;
20'b00011100010011101011: color_data = 12'b000000001111;
20'b00011100010100000101: color_data = 12'b000001101111;
20'b00011100010100000110: color_data = 12'b000001101111;
20'b00011100010100000111: color_data = 12'b000001101111;
20'b00011100010100001000: color_data = 12'b000001101111;
20'b00011100010100001001: color_data = 12'b000001101111;
20'b00011100010100001010: color_data = 12'b000001101111;
20'b00011100010100001011: color_data = 12'b000001101111;
20'b00011100010100001100: color_data = 12'b000001101111;
20'b00011100010100001101: color_data = 12'b000001101111;
20'b00011100010100001110: color_data = 12'b000001101111;
20'b00011100010100001111: color_data = 12'b000001101111;
20'b00011100010100010000: color_data = 12'b000001101111;
20'b00011100010100010001: color_data = 12'b000001101111;
20'b00011100010100010010: color_data = 12'b000001101111;
20'b00011100010100010011: color_data = 12'b000001101111;
20'b00011100010100010100: color_data = 12'b000001101111;
20'b00011100010100010101: color_data = 12'b000001101111;
20'b00011100010100010110: color_data = 12'b000001101111;
20'b00011100010100010111: color_data = 12'b000001101111;
20'b00011100010100011000: color_data = 12'b000001101111;
20'b00011100010100011001: color_data = 12'b000001101111;
20'b00011100010100011010: color_data = 12'b000001101111;
20'b00011100010100011011: color_data = 12'b000001101111;
20'b00011100010100011100: color_data = 12'b000001101111;
20'b00011100010100011101: color_data = 12'b000001101111;
20'b00011100010100011110: color_data = 12'b000001101111;
20'b00011100010100011111: color_data = 12'b000001101111;
20'b00011100010100100000: color_data = 12'b000001101111;
20'b00011100010100100001: color_data = 12'b000001101111;
20'b00011100010100100010: color_data = 12'b000001101111;
20'b00011100010100100011: color_data = 12'b000001101111;
20'b00011100010100100100: color_data = 12'b000001101111;
20'b00011100010100111110: color_data = 12'b000011111111;
20'b00011100010100111111: color_data = 12'b000011111111;
20'b00011100010101000000: color_data = 12'b000011111111;
20'b00011100010101000001: color_data = 12'b000011111111;
20'b00011100010101000010: color_data = 12'b000011111111;
20'b00011100010101000011: color_data = 12'b000011111111;
20'b00011100010101000100: color_data = 12'b000011111111;
20'b00011100010101000101: color_data = 12'b000011111111;
20'b00011100010101011111: color_data = 12'b111101110000;
20'b00011100010101100000: color_data = 12'b111101110000;
20'b00011100010101100001: color_data = 12'b111101110000;
20'b00011100010101100010: color_data = 12'b111101110000;
20'b00011100010101100011: color_data = 12'b111101110000;
20'b00011100010101100100: color_data = 12'b111101110000;
20'b00011100010101100101: color_data = 12'b111101110000;
20'b00011100010101100110: color_data = 12'b111101110000;
20'b00011100010101100111: color_data = 12'b111101110000;
20'b00011100010101101000: color_data = 12'b111101110000;
20'b00011100010101101001: color_data = 12'b111101110000;
20'b00011100010101101010: color_data = 12'b111101110000;
20'b00011100010101101011: color_data = 12'b111101110000;
20'b00011100010101101100: color_data = 12'b111101110000;
20'b00011100010101101101: color_data = 12'b111101110000;
20'b00011100010101101110: color_data = 12'b111101110000;
20'b00011100010101101111: color_data = 12'b111101110000;
20'b00011100010101110000: color_data = 12'b111101110000;
20'b00011100010101110001: color_data = 12'b111101110000;
20'b00011100010101110010: color_data = 12'b111101110000;
20'b00011100010101110011: color_data = 12'b111101110000;
20'b00011100010101110100: color_data = 12'b111101110000;
20'b00011100010101110101: color_data = 12'b111101110000;
20'b00011100010101110110: color_data = 12'b111101110000;
20'b00011100010110000111: color_data = 12'b000011110000;
20'b00011100010110001000: color_data = 12'b000011110000;
20'b00011100010110001001: color_data = 12'b000011110000;
20'b00011100010110001010: color_data = 12'b000011110000;
20'b00011100010110001011: color_data = 12'b000011110000;
20'b00011100010110001100: color_data = 12'b000011110000;
20'b00011100010110001101: color_data = 12'b000011110000;
20'b00011100010110001110: color_data = 12'b000011110000;
20'b00011100010110001111: color_data = 12'b000011110000;
20'b00011100010110011000: color_data = 12'b111100001111;
20'b00011100010110011001: color_data = 12'b111100001111;
20'b00011100010110011010: color_data = 12'b111100001111;
20'b00011100010110011011: color_data = 12'b111100001111;
20'b00011100010110011100: color_data = 12'b111100001111;
20'b00011100010110011101: color_data = 12'b111100001111;
20'b00011100010110011110: color_data = 12'b111100001111;
20'b00011100010110011111: color_data = 12'b111100001111;
20'b00011100010110100000: color_data = 12'b111100001111;
20'b00011100010110100001: color_data = 12'b111100001111;
20'b00011100010110100010: color_data = 12'b111100001111;
20'b00011100010110100011: color_data = 12'b111100001111;
20'b00011100010110100100: color_data = 12'b111100001111;
20'b00011100010110100101: color_data = 12'b111100001111;
20'b00011100010110100110: color_data = 12'b111100001111;
20'b00011100010110100111: color_data = 12'b111100001111;
20'b00011100010110101000: color_data = 12'b111100001111;
20'b00011100010110101001: color_data = 12'b111100001111;
20'b00011100010110101010: color_data = 12'b111100001111;
20'b00011100010110101011: color_data = 12'b111100001111;
20'b00011100010110101100: color_data = 12'b111100001111;
20'b00011100010110101101: color_data = 12'b111100001111;
20'b00011100010110101110: color_data = 12'b111100001111;
20'b00011100010110101111: color_data = 12'b111100001111;
20'b00011100010110110000: color_data = 12'b111100001111;
20'b00011100010110110001: color_data = 12'b111100001111;
20'b00011100010110110010: color_data = 12'b111100001111;
20'b00011100010110110011: color_data = 12'b111100001111;
20'b00011100010110110100: color_data = 12'b111100001111;
20'b00011100010110110101: color_data = 12'b111100001111;
20'b00011100010110110110: color_data = 12'b111100001111;
20'b00011100010110110111: color_data = 12'b111100001111;
20'b00011100100011100100: color_data = 12'b000000001111;
20'b00011100100011100101: color_data = 12'b000000001111;
20'b00011100100011100110: color_data = 12'b000000001111;
20'b00011100100011100111: color_data = 12'b000000001111;
20'b00011100100011101000: color_data = 12'b000000001111;
20'b00011100100011101001: color_data = 12'b000000001111;
20'b00011100100011101010: color_data = 12'b000000001111;
20'b00011100100011101011: color_data = 12'b000000001111;
20'b00011100100100000101: color_data = 12'b000001101111;
20'b00011100100100000110: color_data = 12'b000001101111;
20'b00011100100100000111: color_data = 12'b000001101111;
20'b00011100100100001000: color_data = 12'b000001101111;
20'b00011100100100001001: color_data = 12'b000001101111;
20'b00011100100100001010: color_data = 12'b000001101111;
20'b00011100100100001011: color_data = 12'b000001101111;
20'b00011100100100001100: color_data = 12'b000001101111;
20'b00011100100100001101: color_data = 12'b000001101111;
20'b00011100100100001110: color_data = 12'b000001101111;
20'b00011100100100001111: color_data = 12'b000001101111;
20'b00011100100100010000: color_data = 12'b000001101111;
20'b00011100100100010001: color_data = 12'b000001101111;
20'b00011100100100010010: color_data = 12'b000001101111;
20'b00011100100100010011: color_data = 12'b000001101111;
20'b00011100100100010100: color_data = 12'b000001101111;
20'b00011100100100010101: color_data = 12'b000001101111;
20'b00011100100100010110: color_data = 12'b000001101111;
20'b00011100100100010111: color_data = 12'b000001101111;
20'b00011100100100011000: color_data = 12'b000001101111;
20'b00011100100100011001: color_data = 12'b000001101111;
20'b00011100100100011010: color_data = 12'b000001101111;
20'b00011100100100011011: color_data = 12'b000001101111;
20'b00011100100100011100: color_data = 12'b000001101111;
20'b00011100100100011101: color_data = 12'b000001101111;
20'b00011100100100011110: color_data = 12'b000001101111;
20'b00011100100100011111: color_data = 12'b000001101111;
20'b00011100100100100000: color_data = 12'b000001101111;
20'b00011100100100100001: color_data = 12'b000001101111;
20'b00011100100100100010: color_data = 12'b000001101111;
20'b00011100100100100011: color_data = 12'b000001101111;
20'b00011100100100100100: color_data = 12'b000001101111;
20'b00011100100100111110: color_data = 12'b000011111111;
20'b00011100100100111111: color_data = 12'b000011111111;
20'b00011100100101000000: color_data = 12'b000011111111;
20'b00011100100101000001: color_data = 12'b000011111111;
20'b00011100100101000010: color_data = 12'b000011111111;
20'b00011100100101000011: color_data = 12'b000011111111;
20'b00011100100101000100: color_data = 12'b000011111111;
20'b00011100100101000101: color_data = 12'b000011111111;
20'b00011100100101011111: color_data = 12'b111101110000;
20'b00011100100101100000: color_data = 12'b111101110000;
20'b00011100100101100001: color_data = 12'b111101110000;
20'b00011100100101100010: color_data = 12'b111101110000;
20'b00011100100101100011: color_data = 12'b111101110000;
20'b00011100100101100100: color_data = 12'b111101110000;
20'b00011100100101100101: color_data = 12'b111101110000;
20'b00011100100101100110: color_data = 12'b111101110000;
20'b00011100100101100111: color_data = 12'b111101110000;
20'b00011100100101101000: color_data = 12'b111101110000;
20'b00011100100101101001: color_data = 12'b111101110000;
20'b00011100100101101010: color_data = 12'b111101110000;
20'b00011100100101101011: color_data = 12'b111101110000;
20'b00011100100101101100: color_data = 12'b111101110000;
20'b00011100100101101101: color_data = 12'b111101110000;
20'b00011100100101101110: color_data = 12'b111101110000;
20'b00011100100101101111: color_data = 12'b111101110000;
20'b00011100100101110000: color_data = 12'b111101110000;
20'b00011100100101110001: color_data = 12'b111101110000;
20'b00011100100101110010: color_data = 12'b111101110000;
20'b00011100100101110011: color_data = 12'b111101110000;
20'b00011100100101110100: color_data = 12'b111101110000;
20'b00011100100101110101: color_data = 12'b111101110000;
20'b00011100100101110110: color_data = 12'b111101110000;
20'b00011100100110000111: color_data = 12'b000011110000;
20'b00011100100110001000: color_data = 12'b000011110000;
20'b00011100100110001001: color_data = 12'b000011110000;
20'b00011100100110001010: color_data = 12'b000011110000;
20'b00011100100110001011: color_data = 12'b000011110000;
20'b00011100100110001100: color_data = 12'b000011110000;
20'b00011100100110001101: color_data = 12'b000011110000;
20'b00011100100110001110: color_data = 12'b000011110000;
20'b00011100100110001111: color_data = 12'b000011110000;
20'b00011100100110011000: color_data = 12'b111100001111;
20'b00011100100110011001: color_data = 12'b111100001111;
20'b00011100100110011010: color_data = 12'b111100001111;
20'b00011100100110011011: color_data = 12'b111100001111;
20'b00011100100110011100: color_data = 12'b111100001111;
20'b00011100100110011101: color_data = 12'b111100001111;
20'b00011100100110011110: color_data = 12'b111100001111;
20'b00011100100110011111: color_data = 12'b111100001111;
20'b00011100100110100000: color_data = 12'b111100001111;
20'b00011100100110100001: color_data = 12'b111100001111;
20'b00011100100110100010: color_data = 12'b111100001111;
20'b00011100100110100011: color_data = 12'b111100001111;
20'b00011100100110100100: color_data = 12'b111100001111;
20'b00011100100110100101: color_data = 12'b111100001111;
20'b00011100100110100110: color_data = 12'b111100001111;
20'b00011100100110100111: color_data = 12'b111100001111;
20'b00011100100110101000: color_data = 12'b111100001111;
20'b00011100100110101001: color_data = 12'b111100001111;
20'b00011100100110101010: color_data = 12'b111100001111;
20'b00011100100110101011: color_data = 12'b111100001111;
20'b00011100100110101100: color_data = 12'b111100001111;
20'b00011100100110101101: color_data = 12'b111100001111;
20'b00011100100110101110: color_data = 12'b111100001111;
20'b00011100100110101111: color_data = 12'b111100001111;
20'b00011100100110110000: color_data = 12'b111100001111;
20'b00011100100110110001: color_data = 12'b111100001111;
20'b00011100100110110010: color_data = 12'b111100001111;
20'b00011100100110110011: color_data = 12'b111100001111;
20'b00011100100110110100: color_data = 12'b111100001111;
20'b00011100100110110101: color_data = 12'b111100001111;
20'b00011100100110110110: color_data = 12'b111100001111;
20'b00011100100110110111: color_data = 12'b111100001111;
20'b00011100110011100100: color_data = 12'b000000001111;
20'b00011100110011100101: color_data = 12'b000000001111;
20'b00011100110011100110: color_data = 12'b000000001111;
20'b00011100110011100111: color_data = 12'b000000001111;
20'b00011100110011101000: color_data = 12'b000000001111;
20'b00011100110011101001: color_data = 12'b000000001111;
20'b00011100110011101010: color_data = 12'b000000001111;
20'b00011100110011101011: color_data = 12'b000000001111;
20'b00011100110100000101: color_data = 12'b000001101111;
20'b00011100110100000110: color_data = 12'b000001101111;
20'b00011100110100000111: color_data = 12'b000001101111;
20'b00011100110100001000: color_data = 12'b000001101111;
20'b00011100110100001001: color_data = 12'b000001101111;
20'b00011100110100001010: color_data = 12'b000001101111;
20'b00011100110100001011: color_data = 12'b000001101111;
20'b00011100110100001100: color_data = 12'b000001101111;
20'b00011100110100001101: color_data = 12'b000001101111;
20'b00011100110100001110: color_data = 12'b000001101111;
20'b00011100110100001111: color_data = 12'b000001101111;
20'b00011100110100010000: color_data = 12'b000001101111;
20'b00011100110100010001: color_data = 12'b000001101111;
20'b00011100110100010010: color_data = 12'b000001101111;
20'b00011100110100010011: color_data = 12'b000001101111;
20'b00011100110100010100: color_data = 12'b000001101111;
20'b00011100110100010101: color_data = 12'b000001101111;
20'b00011100110100010110: color_data = 12'b000001101111;
20'b00011100110100010111: color_data = 12'b000001101111;
20'b00011100110100011000: color_data = 12'b000001101111;
20'b00011100110100011001: color_data = 12'b000001101111;
20'b00011100110100011010: color_data = 12'b000001101111;
20'b00011100110100011011: color_data = 12'b000001101111;
20'b00011100110100011100: color_data = 12'b000001101111;
20'b00011100110100011101: color_data = 12'b000001101111;
20'b00011100110100011110: color_data = 12'b000001101111;
20'b00011100110100011111: color_data = 12'b000001101111;
20'b00011100110100100000: color_data = 12'b000001101111;
20'b00011100110100100001: color_data = 12'b000001101111;
20'b00011100110100100010: color_data = 12'b000001101111;
20'b00011100110100100011: color_data = 12'b000001101111;
20'b00011100110100100100: color_data = 12'b000001101111;
20'b00011100110100111110: color_data = 12'b000011111111;
20'b00011100110100111111: color_data = 12'b000011111111;
20'b00011100110101000000: color_data = 12'b000011111111;
20'b00011100110101000001: color_data = 12'b000011111111;
20'b00011100110101000010: color_data = 12'b000011111111;
20'b00011100110101000011: color_data = 12'b000011111111;
20'b00011100110101000100: color_data = 12'b000011111111;
20'b00011100110101000101: color_data = 12'b000011111111;
20'b00011100110101011111: color_data = 12'b111101110000;
20'b00011100110101100000: color_data = 12'b111101110000;
20'b00011100110101100001: color_data = 12'b111101110000;
20'b00011100110101100010: color_data = 12'b111101110000;
20'b00011100110101100011: color_data = 12'b111101110000;
20'b00011100110101100100: color_data = 12'b111101110000;
20'b00011100110101100101: color_data = 12'b111101110000;
20'b00011100110101100110: color_data = 12'b111101110000;
20'b00011100110101100111: color_data = 12'b111101110000;
20'b00011100110101101000: color_data = 12'b111101110000;
20'b00011100110101101001: color_data = 12'b111101110000;
20'b00011100110101101010: color_data = 12'b111101110000;
20'b00011100110101101011: color_data = 12'b111101110000;
20'b00011100110101101100: color_data = 12'b111101110000;
20'b00011100110101101101: color_data = 12'b111101110000;
20'b00011100110101101110: color_data = 12'b111101110000;
20'b00011100110101101111: color_data = 12'b111101110000;
20'b00011100110101110000: color_data = 12'b111101110000;
20'b00011100110101110001: color_data = 12'b111101110000;
20'b00011100110101110010: color_data = 12'b111101110000;
20'b00011100110101110011: color_data = 12'b111101110000;
20'b00011100110101110100: color_data = 12'b111101110000;
20'b00011100110101110101: color_data = 12'b111101110000;
20'b00011100110101110110: color_data = 12'b111101110000;
20'b00011100110110000111: color_data = 12'b000011110000;
20'b00011100110110001000: color_data = 12'b000011110000;
20'b00011100110110001001: color_data = 12'b000011110000;
20'b00011100110110001010: color_data = 12'b000011110000;
20'b00011100110110001011: color_data = 12'b000011110000;
20'b00011100110110001100: color_data = 12'b000011110000;
20'b00011100110110001101: color_data = 12'b000011110000;
20'b00011100110110001110: color_data = 12'b000011110000;
20'b00011100110110001111: color_data = 12'b000011110000;
20'b00011100110110011000: color_data = 12'b111100001111;
20'b00011100110110011001: color_data = 12'b111100001111;
20'b00011100110110011010: color_data = 12'b111100001111;
20'b00011100110110011011: color_data = 12'b111100001111;
20'b00011100110110011100: color_data = 12'b111100001111;
20'b00011100110110011101: color_data = 12'b111100001111;
20'b00011100110110011110: color_data = 12'b111100001111;
20'b00011100110110011111: color_data = 12'b111100001111;
20'b00011100110110100000: color_data = 12'b111100001111;
20'b00011100110110100001: color_data = 12'b111100001111;
20'b00011100110110100010: color_data = 12'b111100001111;
20'b00011100110110100011: color_data = 12'b111100001111;
20'b00011100110110100100: color_data = 12'b111100001111;
20'b00011100110110100101: color_data = 12'b111100001111;
20'b00011100110110100110: color_data = 12'b111100001111;
20'b00011100110110100111: color_data = 12'b111100001111;
20'b00011100110110101000: color_data = 12'b111100001111;
20'b00011100110110101001: color_data = 12'b111100001111;
20'b00011100110110101010: color_data = 12'b111100001111;
20'b00011100110110101011: color_data = 12'b111100001111;
20'b00011100110110101100: color_data = 12'b111100001111;
20'b00011100110110101101: color_data = 12'b111100001111;
20'b00011100110110101110: color_data = 12'b111100001111;
20'b00011100110110101111: color_data = 12'b111100001111;
20'b00011100110110110000: color_data = 12'b111100001111;
20'b00011100110110110001: color_data = 12'b111100001111;
20'b00011100110110110010: color_data = 12'b111100001111;
20'b00011100110110110011: color_data = 12'b111100001111;
20'b00011100110110110100: color_data = 12'b111100001111;
20'b00011100110110110101: color_data = 12'b111100001111;
20'b00011100110110110110: color_data = 12'b111100001111;
20'b00011100110110110111: color_data = 12'b111100001111;
20'b00011101000011100100: color_data = 12'b000000001111;
20'b00011101000011100101: color_data = 12'b000000001111;
20'b00011101000011100110: color_data = 12'b000000001111;
20'b00011101000011100111: color_data = 12'b000000001111;
20'b00011101000011101000: color_data = 12'b000000001111;
20'b00011101000011101001: color_data = 12'b000000001111;
20'b00011101000011101010: color_data = 12'b000000001111;
20'b00011101000011101011: color_data = 12'b000000001111;
20'b00011101000100000101: color_data = 12'b000001101111;
20'b00011101000100000110: color_data = 12'b000001101111;
20'b00011101000100000111: color_data = 12'b000001101111;
20'b00011101000100001000: color_data = 12'b000001101111;
20'b00011101000100001001: color_data = 12'b000001101111;
20'b00011101000100001010: color_data = 12'b000001101111;
20'b00011101000100001011: color_data = 12'b000001101111;
20'b00011101000100001100: color_data = 12'b000001101111;
20'b00011101000100111110: color_data = 12'b000011111111;
20'b00011101000100111111: color_data = 12'b000011111111;
20'b00011101000101000000: color_data = 12'b000011111111;
20'b00011101000101000001: color_data = 12'b000011111111;
20'b00011101000101000010: color_data = 12'b000011111111;
20'b00011101000101000011: color_data = 12'b000011111111;
20'b00011101000101000100: color_data = 12'b000011111111;
20'b00011101000101000101: color_data = 12'b000011111111;
20'b00011101000101011111: color_data = 12'b111101110000;
20'b00011101000101100000: color_data = 12'b111101110000;
20'b00011101000101100001: color_data = 12'b111101110000;
20'b00011101000101100010: color_data = 12'b111101110000;
20'b00011101000101100011: color_data = 12'b111101110000;
20'b00011101000101100100: color_data = 12'b111101110000;
20'b00011101000101100101: color_data = 12'b111101110000;
20'b00011101000101100110: color_data = 12'b111101110000;
20'b00011101000101110111: color_data = 12'b111101100000;
20'b00011101000101111000: color_data = 12'b111101100000;
20'b00011101000101111001: color_data = 12'b111101100000;
20'b00011101000101111010: color_data = 12'b111101100000;
20'b00011101000101111011: color_data = 12'b111101100000;
20'b00011101000101111100: color_data = 12'b111101100000;
20'b00011101000101111101: color_data = 12'b111101100000;
20'b00011101000101111110: color_data = 12'b111101100000;
20'b00011101000110000111: color_data = 12'b000011110000;
20'b00011101000110001000: color_data = 12'b000011110000;
20'b00011101000110001001: color_data = 12'b000011110000;
20'b00011101000110001010: color_data = 12'b000011110000;
20'b00011101000110001011: color_data = 12'b000011110000;
20'b00011101000110001100: color_data = 12'b000011110000;
20'b00011101000110001101: color_data = 12'b000011110000;
20'b00011101000110001110: color_data = 12'b000011110000;
20'b00011101000110001111: color_data = 12'b000011110000;
20'b00011101000110110000: color_data = 12'b111100001111;
20'b00011101000110110001: color_data = 12'b111100001111;
20'b00011101000110110010: color_data = 12'b111100001111;
20'b00011101000110110011: color_data = 12'b111100001111;
20'b00011101000110110100: color_data = 12'b111100001111;
20'b00011101000110110101: color_data = 12'b111100001111;
20'b00011101000110110110: color_data = 12'b111100001111;
20'b00011101000110110111: color_data = 12'b111100001111;
20'b00011101010011100100: color_data = 12'b000000001111;
20'b00011101010011100101: color_data = 12'b000000001111;
20'b00011101010011100110: color_data = 12'b000000001111;
20'b00011101010011100111: color_data = 12'b000000001111;
20'b00011101010011101000: color_data = 12'b000000001111;
20'b00011101010011101001: color_data = 12'b000000001111;
20'b00011101010011101010: color_data = 12'b000000001111;
20'b00011101010011101011: color_data = 12'b000000001111;
20'b00011101010100000101: color_data = 12'b000001101111;
20'b00011101010100000110: color_data = 12'b000001101111;
20'b00011101010100000111: color_data = 12'b000001101111;
20'b00011101010100001000: color_data = 12'b000001101111;
20'b00011101010100001001: color_data = 12'b000001101111;
20'b00011101010100001010: color_data = 12'b000001101111;
20'b00011101010100001011: color_data = 12'b000001101111;
20'b00011101010100001100: color_data = 12'b000001101111;
20'b00011101010100111110: color_data = 12'b000011111111;
20'b00011101010100111111: color_data = 12'b000011111111;
20'b00011101010101000000: color_data = 12'b000011111111;
20'b00011101010101000001: color_data = 12'b000011111111;
20'b00011101010101000010: color_data = 12'b000011111111;
20'b00011101010101000011: color_data = 12'b000011111111;
20'b00011101010101000100: color_data = 12'b000011111111;
20'b00011101010101000101: color_data = 12'b000011111111;
20'b00011101010101011111: color_data = 12'b111101110000;
20'b00011101010101100000: color_data = 12'b111101110000;
20'b00011101010101100001: color_data = 12'b111101110000;
20'b00011101010101100010: color_data = 12'b111101110000;
20'b00011101010101100011: color_data = 12'b111101110000;
20'b00011101010101100100: color_data = 12'b111101110000;
20'b00011101010101100101: color_data = 12'b111101110000;
20'b00011101010101100110: color_data = 12'b111101110000;
20'b00011101010101110111: color_data = 12'b111101100000;
20'b00011101010101111000: color_data = 12'b111101100000;
20'b00011101010101111001: color_data = 12'b111101100000;
20'b00011101010101111010: color_data = 12'b111101100000;
20'b00011101010101111011: color_data = 12'b111101100000;
20'b00011101010101111100: color_data = 12'b111101100000;
20'b00011101010101111101: color_data = 12'b111101100000;
20'b00011101010101111110: color_data = 12'b111101100000;
20'b00011101010110000111: color_data = 12'b000011110000;
20'b00011101010110001000: color_data = 12'b000011110000;
20'b00011101010110001001: color_data = 12'b000011110000;
20'b00011101010110001010: color_data = 12'b000011110000;
20'b00011101010110001011: color_data = 12'b000011110000;
20'b00011101010110001100: color_data = 12'b000011110000;
20'b00011101010110001101: color_data = 12'b000011110000;
20'b00011101010110001110: color_data = 12'b000011110000;
20'b00011101010110001111: color_data = 12'b000011110000;
20'b00011101010110110000: color_data = 12'b111100001111;
20'b00011101010110110001: color_data = 12'b111100001111;
20'b00011101010110110010: color_data = 12'b111100001111;
20'b00011101010110110011: color_data = 12'b111100001111;
20'b00011101010110110100: color_data = 12'b111100001111;
20'b00011101010110110101: color_data = 12'b111100001111;
20'b00011101010110110110: color_data = 12'b111100001111;
20'b00011101010110110111: color_data = 12'b111100001111;
20'b00011101100011100100: color_data = 12'b000000001111;
20'b00011101100011100101: color_data = 12'b000000001111;
20'b00011101100011100110: color_data = 12'b000000001111;
20'b00011101100011100111: color_data = 12'b000000001111;
20'b00011101100011101000: color_data = 12'b000000001111;
20'b00011101100011101001: color_data = 12'b000000001111;
20'b00011101100011101010: color_data = 12'b000000001111;
20'b00011101100011101011: color_data = 12'b000000001111;
20'b00011101100100000101: color_data = 12'b000001101111;
20'b00011101100100000110: color_data = 12'b000001101111;
20'b00011101100100000111: color_data = 12'b000001101111;
20'b00011101100100001000: color_data = 12'b000001101111;
20'b00011101100100001001: color_data = 12'b000001101111;
20'b00011101100100001010: color_data = 12'b000001101111;
20'b00011101100100001011: color_data = 12'b000001101111;
20'b00011101100100001100: color_data = 12'b000001101111;
20'b00011101100100111110: color_data = 12'b000011111111;
20'b00011101100100111111: color_data = 12'b000011111111;
20'b00011101100101000000: color_data = 12'b000011111111;
20'b00011101100101000001: color_data = 12'b000011111111;
20'b00011101100101000010: color_data = 12'b000011111111;
20'b00011101100101000011: color_data = 12'b000011111111;
20'b00011101100101000100: color_data = 12'b000011111111;
20'b00011101100101000101: color_data = 12'b000011111111;
20'b00011101100101011111: color_data = 12'b111101110000;
20'b00011101100101100000: color_data = 12'b111101110000;
20'b00011101100101100001: color_data = 12'b111101110000;
20'b00011101100101100010: color_data = 12'b111101110000;
20'b00011101100101100011: color_data = 12'b111101110000;
20'b00011101100101100100: color_data = 12'b111101110000;
20'b00011101100101100101: color_data = 12'b111101110000;
20'b00011101100101100110: color_data = 12'b111101110000;
20'b00011101100101110111: color_data = 12'b111101100000;
20'b00011101100101111000: color_data = 12'b111101100000;
20'b00011101100101111001: color_data = 12'b111101100000;
20'b00011101100101111010: color_data = 12'b111101100000;
20'b00011101100101111011: color_data = 12'b111101100000;
20'b00011101100101111100: color_data = 12'b111101100000;
20'b00011101100101111101: color_data = 12'b111101100000;
20'b00011101100101111110: color_data = 12'b111101100000;
20'b00011101100110000111: color_data = 12'b000011110000;
20'b00011101100110001000: color_data = 12'b000011110000;
20'b00011101100110001001: color_data = 12'b000011110000;
20'b00011101100110001010: color_data = 12'b000011110000;
20'b00011101100110001011: color_data = 12'b000011110000;
20'b00011101100110001100: color_data = 12'b000011110000;
20'b00011101100110001101: color_data = 12'b000011110000;
20'b00011101100110001110: color_data = 12'b000011110000;
20'b00011101100110001111: color_data = 12'b000011110000;
20'b00011101100110110000: color_data = 12'b111100001111;
20'b00011101100110110001: color_data = 12'b111100001111;
20'b00011101100110110010: color_data = 12'b111100001111;
20'b00011101100110110011: color_data = 12'b111100001111;
20'b00011101100110110100: color_data = 12'b111100001111;
20'b00011101100110110101: color_data = 12'b111100001111;
20'b00011101100110110110: color_data = 12'b111100001111;
20'b00011101100110110111: color_data = 12'b111100001111;
20'b00011101110011100100: color_data = 12'b000000001111;
20'b00011101110011100101: color_data = 12'b000000001111;
20'b00011101110011100110: color_data = 12'b000000001111;
20'b00011101110011100111: color_data = 12'b000000001111;
20'b00011101110011101000: color_data = 12'b000000001111;
20'b00011101110011101001: color_data = 12'b000000001111;
20'b00011101110011101010: color_data = 12'b000000001111;
20'b00011101110011101011: color_data = 12'b000000001111;
20'b00011101110100000101: color_data = 12'b000001101111;
20'b00011101110100000110: color_data = 12'b000001101111;
20'b00011101110100000111: color_data = 12'b000001101111;
20'b00011101110100001000: color_data = 12'b000001101111;
20'b00011101110100001001: color_data = 12'b000001101111;
20'b00011101110100001010: color_data = 12'b000001101111;
20'b00011101110100001011: color_data = 12'b000001101111;
20'b00011101110100001100: color_data = 12'b000001101111;
20'b00011101110100111110: color_data = 12'b000011111111;
20'b00011101110100111111: color_data = 12'b000011111111;
20'b00011101110101000000: color_data = 12'b000011111111;
20'b00011101110101000001: color_data = 12'b000011111111;
20'b00011101110101000010: color_data = 12'b000011111111;
20'b00011101110101000011: color_data = 12'b000011111111;
20'b00011101110101000100: color_data = 12'b000011111111;
20'b00011101110101000101: color_data = 12'b000011111111;
20'b00011101110101011111: color_data = 12'b111101110000;
20'b00011101110101100000: color_data = 12'b111101110000;
20'b00011101110101100001: color_data = 12'b111101110000;
20'b00011101110101100010: color_data = 12'b111101110000;
20'b00011101110101100011: color_data = 12'b111101110000;
20'b00011101110101100100: color_data = 12'b111101110000;
20'b00011101110101100101: color_data = 12'b111101110000;
20'b00011101110101100110: color_data = 12'b111101110000;
20'b00011101110101110111: color_data = 12'b111101100000;
20'b00011101110101111000: color_data = 12'b111101100000;
20'b00011101110101111001: color_data = 12'b111101100000;
20'b00011101110101111010: color_data = 12'b111101100000;
20'b00011101110101111011: color_data = 12'b111101100000;
20'b00011101110101111100: color_data = 12'b111101100000;
20'b00011101110101111101: color_data = 12'b111101100000;
20'b00011101110101111110: color_data = 12'b111101100000;
20'b00011101110110000111: color_data = 12'b000011110000;
20'b00011101110110001000: color_data = 12'b000011110000;
20'b00011101110110001001: color_data = 12'b000011110000;
20'b00011101110110001010: color_data = 12'b000011110000;
20'b00011101110110001011: color_data = 12'b000011110000;
20'b00011101110110001100: color_data = 12'b000011110000;
20'b00011101110110001101: color_data = 12'b000011110000;
20'b00011101110110001110: color_data = 12'b000011110000;
20'b00011101110110001111: color_data = 12'b000011110000;
20'b00011101110110110000: color_data = 12'b111100001111;
20'b00011101110110110001: color_data = 12'b111100001111;
20'b00011101110110110010: color_data = 12'b111100001111;
20'b00011101110110110011: color_data = 12'b111100001111;
20'b00011101110110110100: color_data = 12'b111100001111;
20'b00011101110110110101: color_data = 12'b111100001111;
20'b00011101110110110110: color_data = 12'b111100001111;
20'b00011101110110110111: color_data = 12'b111100001111;
20'b00011110000011100100: color_data = 12'b000000001111;
20'b00011110000011100101: color_data = 12'b000000001111;
20'b00011110000011100110: color_data = 12'b000000001111;
20'b00011110000011100111: color_data = 12'b000000001111;
20'b00011110000011101000: color_data = 12'b000000001111;
20'b00011110000011101001: color_data = 12'b000000001111;
20'b00011110000011101010: color_data = 12'b000000001111;
20'b00011110000011101011: color_data = 12'b000000001111;
20'b00011110000100000101: color_data = 12'b000001101111;
20'b00011110000100000110: color_data = 12'b000001101111;
20'b00011110000100000111: color_data = 12'b000001101111;
20'b00011110000100001000: color_data = 12'b000001101111;
20'b00011110000100001001: color_data = 12'b000001101111;
20'b00011110000100001010: color_data = 12'b000001101111;
20'b00011110000100001011: color_data = 12'b000001101111;
20'b00011110000100001100: color_data = 12'b000001101111;
20'b00011110000100111110: color_data = 12'b000011111111;
20'b00011110000100111111: color_data = 12'b000011111111;
20'b00011110000101000000: color_data = 12'b000011111111;
20'b00011110000101000001: color_data = 12'b000011111111;
20'b00011110000101000010: color_data = 12'b000011111111;
20'b00011110000101000011: color_data = 12'b000011111111;
20'b00011110000101000100: color_data = 12'b000011111111;
20'b00011110000101000101: color_data = 12'b000011111111;
20'b00011110000101011111: color_data = 12'b111101110000;
20'b00011110000101100000: color_data = 12'b111101110000;
20'b00011110000101100001: color_data = 12'b111101110000;
20'b00011110000101100010: color_data = 12'b111101110000;
20'b00011110000101100011: color_data = 12'b111101110000;
20'b00011110000101100100: color_data = 12'b111101110000;
20'b00011110000101100101: color_data = 12'b111101110000;
20'b00011110000101100110: color_data = 12'b111101110000;
20'b00011110000101110111: color_data = 12'b111101100000;
20'b00011110000101111000: color_data = 12'b111101100000;
20'b00011110000101111001: color_data = 12'b111101100000;
20'b00011110000101111010: color_data = 12'b111101100000;
20'b00011110000101111011: color_data = 12'b111101100000;
20'b00011110000101111100: color_data = 12'b111101100000;
20'b00011110000101111101: color_data = 12'b111101100000;
20'b00011110000101111110: color_data = 12'b111101100000;
20'b00011110000110000111: color_data = 12'b000011110000;
20'b00011110000110001000: color_data = 12'b000011110000;
20'b00011110000110001001: color_data = 12'b000011110000;
20'b00011110000110001010: color_data = 12'b000011110000;
20'b00011110000110001011: color_data = 12'b000011110000;
20'b00011110000110001100: color_data = 12'b000011110000;
20'b00011110000110001101: color_data = 12'b000011110000;
20'b00011110000110001110: color_data = 12'b000011110000;
20'b00011110000110001111: color_data = 12'b000011110000;
20'b00011110000110110000: color_data = 12'b111100001111;
20'b00011110000110110001: color_data = 12'b111100001111;
20'b00011110000110110010: color_data = 12'b111100001111;
20'b00011110000110110011: color_data = 12'b111100001111;
20'b00011110000110110100: color_data = 12'b111100001111;
20'b00011110000110110101: color_data = 12'b111100001111;
20'b00011110000110110110: color_data = 12'b111100001111;
20'b00011110000110110111: color_data = 12'b111100001111;
20'b00011110010011100100: color_data = 12'b000000001111;
20'b00011110010011100101: color_data = 12'b000000001111;
20'b00011110010011100110: color_data = 12'b000000001111;
20'b00011110010011100111: color_data = 12'b000000001111;
20'b00011110010011101000: color_data = 12'b000000001111;
20'b00011110010011101001: color_data = 12'b000000001111;
20'b00011110010011101010: color_data = 12'b000000001111;
20'b00011110010011101011: color_data = 12'b000000001111;
20'b00011110010100000101: color_data = 12'b000001101111;
20'b00011110010100000110: color_data = 12'b000001101111;
20'b00011110010100000111: color_data = 12'b000001101111;
20'b00011110010100001000: color_data = 12'b000001101111;
20'b00011110010100001001: color_data = 12'b000001101111;
20'b00011110010100001010: color_data = 12'b000001101111;
20'b00011110010100001011: color_data = 12'b000001101111;
20'b00011110010100001100: color_data = 12'b000001101111;
20'b00011110010100111110: color_data = 12'b000011111111;
20'b00011110010100111111: color_data = 12'b000011111111;
20'b00011110010101000000: color_data = 12'b000011111111;
20'b00011110010101000001: color_data = 12'b000011111111;
20'b00011110010101000010: color_data = 12'b000011111111;
20'b00011110010101000011: color_data = 12'b000011111111;
20'b00011110010101000100: color_data = 12'b000011111111;
20'b00011110010101000101: color_data = 12'b000011111111;
20'b00011110010101011111: color_data = 12'b111101110000;
20'b00011110010101100000: color_data = 12'b111101110000;
20'b00011110010101100001: color_data = 12'b111101110000;
20'b00011110010101100010: color_data = 12'b111101110000;
20'b00011110010101100011: color_data = 12'b111101110000;
20'b00011110010101100100: color_data = 12'b111101110000;
20'b00011110010101100101: color_data = 12'b111101110000;
20'b00011110010101100110: color_data = 12'b111101110000;
20'b00011110010101110111: color_data = 12'b111101100000;
20'b00011110010101111000: color_data = 12'b111101100000;
20'b00011110010101111001: color_data = 12'b111101100000;
20'b00011110010101111010: color_data = 12'b111101100000;
20'b00011110010101111011: color_data = 12'b111101100000;
20'b00011110010101111100: color_data = 12'b111101100000;
20'b00011110010101111101: color_data = 12'b111101100000;
20'b00011110010101111110: color_data = 12'b111101100000;
20'b00011110010110000111: color_data = 12'b000011110000;
20'b00011110010110001000: color_data = 12'b000011110000;
20'b00011110010110001001: color_data = 12'b000011110000;
20'b00011110010110001010: color_data = 12'b000011110000;
20'b00011110010110001011: color_data = 12'b000011110000;
20'b00011110010110001100: color_data = 12'b000011110000;
20'b00011110010110001101: color_data = 12'b000011110000;
20'b00011110010110001110: color_data = 12'b000011110000;
20'b00011110010110001111: color_data = 12'b000011110000;
20'b00011110010110110000: color_data = 12'b111100001111;
20'b00011110010110110001: color_data = 12'b111100001111;
20'b00011110010110110010: color_data = 12'b111100001111;
20'b00011110010110110011: color_data = 12'b111100001111;
20'b00011110010110110100: color_data = 12'b111100001111;
20'b00011110010110110101: color_data = 12'b111100001111;
20'b00011110010110110110: color_data = 12'b111100001111;
20'b00011110010110110111: color_data = 12'b111100001111;
20'b00011110100011100100: color_data = 12'b000000001111;
20'b00011110100011100101: color_data = 12'b000000001111;
20'b00011110100011100110: color_data = 12'b000000001111;
20'b00011110100011100111: color_data = 12'b000000001111;
20'b00011110100011101000: color_data = 12'b000000001111;
20'b00011110100011101001: color_data = 12'b000000001111;
20'b00011110100011101010: color_data = 12'b000000001111;
20'b00011110100011101011: color_data = 12'b000000001111;
20'b00011110100100000101: color_data = 12'b000001101111;
20'b00011110100100000110: color_data = 12'b000001101111;
20'b00011110100100000111: color_data = 12'b000001101111;
20'b00011110100100001000: color_data = 12'b000001101111;
20'b00011110100100001001: color_data = 12'b000001101111;
20'b00011110100100001010: color_data = 12'b000001101111;
20'b00011110100100001011: color_data = 12'b000001101111;
20'b00011110100100001100: color_data = 12'b000001101111;
20'b00011110100100111110: color_data = 12'b000011111111;
20'b00011110100100111111: color_data = 12'b000011111111;
20'b00011110100101000000: color_data = 12'b000011111111;
20'b00011110100101000001: color_data = 12'b000011111111;
20'b00011110100101000010: color_data = 12'b000011111111;
20'b00011110100101000011: color_data = 12'b000011111111;
20'b00011110100101000100: color_data = 12'b000011111111;
20'b00011110100101000101: color_data = 12'b000011111111;
20'b00011110100101011111: color_data = 12'b111101110000;
20'b00011110100101100000: color_data = 12'b111101110000;
20'b00011110100101100001: color_data = 12'b111101110000;
20'b00011110100101100010: color_data = 12'b111101110000;
20'b00011110100101100011: color_data = 12'b111101110000;
20'b00011110100101100100: color_data = 12'b111101110000;
20'b00011110100101100101: color_data = 12'b111101110000;
20'b00011110100101100110: color_data = 12'b111101110000;
20'b00011110100101110111: color_data = 12'b111101100000;
20'b00011110100101111000: color_data = 12'b111101100000;
20'b00011110100101111001: color_data = 12'b111101100000;
20'b00011110100101111010: color_data = 12'b111101100000;
20'b00011110100101111011: color_data = 12'b111101100000;
20'b00011110100101111100: color_data = 12'b111101100000;
20'b00011110100101111101: color_data = 12'b111101100000;
20'b00011110100101111110: color_data = 12'b111101100000;
20'b00011110100110000111: color_data = 12'b000011110000;
20'b00011110100110001000: color_data = 12'b000011110000;
20'b00011110100110001001: color_data = 12'b000011110000;
20'b00011110100110001010: color_data = 12'b000011110000;
20'b00011110100110001011: color_data = 12'b000011110000;
20'b00011110100110001100: color_data = 12'b000011110000;
20'b00011110100110001101: color_data = 12'b000011110000;
20'b00011110100110001110: color_data = 12'b000011110000;
20'b00011110100110001111: color_data = 12'b000011110000;
20'b00011110100110110000: color_data = 12'b111100001111;
20'b00011110100110110001: color_data = 12'b111100001111;
20'b00011110100110110010: color_data = 12'b111100001111;
20'b00011110100110110011: color_data = 12'b111100001111;
20'b00011110100110110100: color_data = 12'b111100001111;
20'b00011110100110110101: color_data = 12'b111100001111;
20'b00011110100110110110: color_data = 12'b111100001111;
20'b00011110100110110111: color_data = 12'b111100001111;
20'b00011110110011100100: color_data = 12'b000000001111;
20'b00011110110011100101: color_data = 12'b000000001111;
20'b00011110110011100110: color_data = 12'b000000001111;
20'b00011110110011100111: color_data = 12'b000000001111;
20'b00011110110011101000: color_data = 12'b000000001111;
20'b00011110110011101001: color_data = 12'b000000001111;
20'b00011110110011101010: color_data = 12'b000000001111;
20'b00011110110011101011: color_data = 12'b000000001111;
20'b00011110110100000101: color_data = 12'b000001101111;
20'b00011110110100000110: color_data = 12'b000001101111;
20'b00011110110100000111: color_data = 12'b000001101111;
20'b00011110110100001000: color_data = 12'b000001101111;
20'b00011110110100001001: color_data = 12'b000001101111;
20'b00011110110100001010: color_data = 12'b000001101111;
20'b00011110110100001011: color_data = 12'b000001101111;
20'b00011110110100001100: color_data = 12'b000001101111;
20'b00011110110100111110: color_data = 12'b000011111111;
20'b00011110110100111111: color_data = 12'b000011111111;
20'b00011110110101000000: color_data = 12'b000011111111;
20'b00011110110101000001: color_data = 12'b000011111111;
20'b00011110110101000010: color_data = 12'b000011111111;
20'b00011110110101000011: color_data = 12'b000011111111;
20'b00011110110101000100: color_data = 12'b000011111111;
20'b00011110110101000101: color_data = 12'b000011111111;
20'b00011110110101011111: color_data = 12'b111101110000;
20'b00011110110101100000: color_data = 12'b111101110000;
20'b00011110110101100001: color_data = 12'b111101110000;
20'b00011110110101100010: color_data = 12'b111101110000;
20'b00011110110101100011: color_data = 12'b111101110000;
20'b00011110110101100100: color_data = 12'b111101110000;
20'b00011110110101100101: color_data = 12'b111101110000;
20'b00011110110101100110: color_data = 12'b111101110000;
20'b00011110110101110111: color_data = 12'b111101100000;
20'b00011110110101111000: color_data = 12'b111101100000;
20'b00011110110101111001: color_data = 12'b111101100000;
20'b00011110110101111010: color_data = 12'b111101100000;
20'b00011110110101111011: color_data = 12'b111101100000;
20'b00011110110101111100: color_data = 12'b111101100000;
20'b00011110110101111101: color_data = 12'b111101100000;
20'b00011110110101111110: color_data = 12'b111101100000;
20'b00011110110110000111: color_data = 12'b000011110000;
20'b00011110110110001000: color_data = 12'b000011110000;
20'b00011110110110001001: color_data = 12'b000011110000;
20'b00011110110110001010: color_data = 12'b000011110000;
20'b00011110110110001011: color_data = 12'b000011110000;
20'b00011110110110001100: color_data = 12'b000011110000;
20'b00011110110110001101: color_data = 12'b000011110000;
20'b00011110110110001110: color_data = 12'b000011110000;
20'b00011110110110001111: color_data = 12'b000011110000;
20'b00011110110110110000: color_data = 12'b111100001111;
20'b00011110110110110001: color_data = 12'b111100001111;
20'b00011110110110110010: color_data = 12'b111100001111;
20'b00011110110110110011: color_data = 12'b111100001111;
20'b00011110110110110100: color_data = 12'b111100001111;
20'b00011110110110110101: color_data = 12'b111100001111;
20'b00011110110110110110: color_data = 12'b111100001111;
20'b00011110110110110111: color_data = 12'b111100001111;
20'b00011111000011100100: color_data = 12'b000000001111;
20'b00011111000011100101: color_data = 12'b000000001111;
20'b00011111000011100110: color_data = 12'b000000001111;
20'b00011111000011100111: color_data = 12'b000000001111;
20'b00011111000011101000: color_data = 12'b000000001111;
20'b00011111000011101001: color_data = 12'b000000001111;
20'b00011111000011101010: color_data = 12'b000000001111;
20'b00011111000011101011: color_data = 12'b000000001111;
20'b00011111000100000101: color_data = 12'b000001101111;
20'b00011111000100000110: color_data = 12'b000001101111;
20'b00011111000100000111: color_data = 12'b000001101111;
20'b00011111000100001000: color_data = 12'b000001101111;
20'b00011111000100001001: color_data = 12'b000001101111;
20'b00011111000100001010: color_data = 12'b000001101111;
20'b00011111000100001011: color_data = 12'b000001101111;
20'b00011111000100001100: color_data = 12'b000001101111;
20'b00011111000100111110: color_data = 12'b000011111111;
20'b00011111000100111111: color_data = 12'b000011111111;
20'b00011111000101000000: color_data = 12'b000011111111;
20'b00011111000101000001: color_data = 12'b000011111111;
20'b00011111000101000010: color_data = 12'b000011111111;
20'b00011111000101000011: color_data = 12'b000011111111;
20'b00011111000101000100: color_data = 12'b000011111111;
20'b00011111000101000101: color_data = 12'b000011111111;
20'b00011111000101011111: color_data = 12'b111101110000;
20'b00011111000101100000: color_data = 12'b111101110000;
20'b00011111000101100001: color_data = 12'b111101110000;
20'b00011111000101100010: color_data = 12'b111101110000;
20'b00011111000101100011: color_data = 12'b111101110000;
20'b00011111000101100100: color_data = 12'b111101110000;
20'b00011111000101100101: color_data = 12'b111101110000;
20'b00011111000101100110: color_data = 12'b111101110000;
20'b00011111000101110111: color_data = 12'b111101100000;
20'b00011111000101111000: color_data = 12'b111101100000;
20'b00011111000101111001: color_data = 12'b111101100000;
20'b00011111000101111010: color_data = 12'b111101100000;
20'b00011111000101111011: color_data = 12'b111101100000;
20'b00011111000101111100: color_data = 12'b111101100000;
20'b00011111000101111101: color_data = 12'b111101100000;
20'b00011111000101111110: color_data = 12'b111101100000;
20'b00011111000110000111: color_data = 12'b000011110000;
20'b00011111000110001000: color_data = 12'b000011110000;
20'b00011111000110001001: color_data = 12'b000011110000;
20'b00011111000110001010: color_data = 12'b000011110000;
20'b00011111000110001011: color_data = 12'b000011110000;
20'b00011111000110001100: color_data = 12'b000011110000;
20'b00011111000110001101: color_data = 12'b000011110000;
20'b00011111000110001110: color_data = 12'b000011110000;
20'b00011111000110001111: color_data = 12'b000011110000;
20'b00011111000110110000: color_data = 12'b111100001111;
20'b00011111000110110001: color_data = 12'b111100001111;
20'b00011111000110110010: color_data = 12'b111100001111;
20'b00011111000110110011: color_data = 12'b111100001111;
20'b00011111000110110100: color_data = 12'b111100001111;
20'b00011111000110110101: color_data = 12'b111100001111;
20'b00011111000110110110: color_data = 12'b111100001111;
20'b00011111000110110111: color_data = 12'b111100001111;
20'b00011111010011100100: color_data = 12'b000000001111;
20'b00011111010011100101: color_data = 12'b000000001111;
20'b00011111010011100110: color_data = 12'b000000001111;
20'b00011111010011100111: color_data = 12'b000000001111;
20'b00011111010011101000: color_data = 12'b000000001111;
20'b00011111010011101001: color_data = 12'b000000001111;
20'b00011111010011101010: color_data = 12'b000000001111;
20'b00011111010011101011: color_data = 12'b000000001111;
20'b00011111010100000101: color_data = 12'b000001101111;
20'b00011111010100000110: color_data = 12'b000001101111;
20'b00011111010100000111: color_data = 12'b000001101111;
20'b00011111010100001000: color_data = 12'b000001101111;
20'b00011111010100001001: color_data = 12'b000001101111;
20'b00011111010100001010: color_data = 12'b000001101111;
20'b00011111010100001011: color_data = 12'b000001101111;
20'b00011111010100001100: color_data = 12'b000001101111;
20'b00011111010100111110: color_data = 12'b000011111111;
20'b00011111010100111111: color_data = 12'b000011111111;
20'b00011111010101000000: color_data = 12'b000011111111;
20'b00011111010101000001: color_data = 12'b000011111111;
20'b00011111010101000010: color_data = 12'b000011111111;
20'b00011111010101000011: color_data = 12'b000011111111;
20'b00011111010101000100: color_data = 12'b000011111111;
20'b00011111010101000101: color_data = 12'b000011111111;
20'b00011111010101011111: color_data = 12'b111101110000;
20'b00011111010101100000: color_data = 12'b111101110000;
20'b00011111010101100001: color_data = 12'b111101110000;
20'b00011111010101100010: color_data = 12'b111101110000;
20'b00011111010101100011: color_data = 12'b111101110000;
20'b00011111010101100100: color_data = 12'b111101110000;
20'b00011111010101100101: color_data = 12'b111101110000;
20'b00011111010101100110: color_data = 12'b111101110000;
20'b00011111010101110111: color_data = 12'b111101100000;
20'b00011111010101111000: color_data = 12'b111101100000;
20'b00011111010101111001: color_data = 12'b111101100000;
20'b00011111010101111010: color_data = 12'b111101100000;
20'b00011111010101111011: color_data = 12'b111101100000;
20'b00011111010101111100: color_data = 12'b111101100000;
20'b00011111010101111101: color_data = 12'b111101100000;
20'b00011111010101111110: color_data = 12'b111101100000;
20'b00011111010110000111: color_data = 12'b000011110000;
20'b00011111010110001000: color_data = 12'b000011110000;
20'b00011111010110001001: color_data = 12'b000011110000;
20'b00011111010110001010: color_data = 12'b000011110000;
20'b00011111010110001011: color_data = 12'b000011110000;
20'b00011111010110001100: color_data = 12'b000011110000;
20'b00011111010110001101: color_data = 12'b000011110000;
20'b00011111010110001110: color_data = 12'b000011110000;
20'b00011111010110001111: color_data = 12'b000011110000;
20'b00011111010110110000: color_data = 12'b111100001111;
20'b00011111010110110001: color_data = 12'b111100001111;
20'b00011111010110110010: color_data = 12'b111100001111;
20'b00011111010110110011: color_data = 12'b111100001111;
20'b00011111010110110100: color_data = 12'b111100001111;
20'b00011111010110110101: color_data = 12'b111100001111;
20'b00011111010110110110: color_data = 12'b111100001111;
20'b00011111010110110111: color_data = 12'b111100001111;
20'b00011111100011100100: color_data = 12'b000000001111;
20'b00011111100011100101: color_data = 12'b000000001111;
20'b00011111100011100110: color_data = 12'b000000001111;
20'b00011111100011100111: color_data = 12'b000000001111;
20'b00011111100011101000: color_data = 12'b000000001111;
20'b00011111100011101001: color_data = 12'b000000001111;
20'b00011111100011101010: color_data = 12'b000000001111;
20'b00011111100011101011: color_data = 12'b000000001111;
20'b00011111100100000101: color_data = 12'b000001101111;
20'b00011111100100000110: color_data = 12'b000001101111;
20'b00011111100100000111: color_data = 12'b000001101111;
20'b00011111100100001000: color_data = 12'b000001101111;
20'b00011111100100001001: color_data = 12'b000001101111;
20'b00011111100100001010: color_data = 12'b000001101111;
20'b00011111100100001011: color_data = 12'b000001101111;
20'b00011111100100001100: color_data = 12'b000001101111;
20'b00011111100100111110: color_data = 12'b000011111111;
20'b00011111100100111111: color_data = 12'b000011111111;
20'b00011111100101000000: color_data = 12'b000011111111;
20'b00011111100101000001: color_data = 12'b000011111111;
20'b00011111100101000010: color_data = 12'b000011111111;
20'b00011111100101000011: color_data = 12'b000011111111;
20'b00011111100101000100: color_data = 12'b000011111111;
20'b00011111100101000101: color_data = 12'b000011111111;
20'b00011111100101011111: color_data = 12'b111101110000;
20'b00011111100101100000: color_data = 12'b111101110000;
20'b00011111100101100001: color_data = 12'b111101110000;
20'b00011111100101100010: color_data = 12'b111101110000;
20'b00011111100101100011: color_data = 12'b111101110000;
20'b00011111100101100100: color_data = 12'b111101110000;
20'b00011111100101100101: color_data = 12'b111101110000;
20'b00011111100101100110: color_data = 12'b111101110000;
20'b00011111100101110111: color_data = 12'b111101100000;
20'b00011111100101111000: color_data = 12'b111101100000;
20'b00011111100101111001: color_data = 12'b111101100000;
20'b00011111100101111010: color_data = 12'b111101100000;
20'b00011111100101111011: color_data = 12'b111101100000;
20'b00011111100101111100: color_data = 12'b111101100000;
20'b00011111100101111101: color_data = 12'b111101100000;
20'b00011111100101111110: color_data = 12'b111101100000;
20'b00011111100110000111: color_data = 12'b000011110000;
20'b00011111100110001000: color_data = 12'b000011110000;
20'b00011111100110001001: color_data = 12'b000011110000;
20'b00011111100110001010: color_data = 12'b000011110000;
20'b00011111100110001011: color_data = 12'b000011110000;
20'b00011111100110001100: color_data = 12'b000011110000;
20'b00011111100110001101: color_data = 12'b000011110000;
20'b00011111100110001110: color_data = 12'b000011110000;
20'b00011111100110001111: color_data = 12'b000011110000;
20'b00011111100110110000: color_data = 12'b111100001111;
20'b00011111100110110001: color_data = 12'b111100001111;
20'b00011111100110110010: color_data = 12'b111100001111;
20'b00011111100110110011: color_data = 12'b111100001111;
20'b00011111100110110100: color_data = 12'b111100001111;
20'b00011111100110110101: color_data = 12'b111100001111;
20'b00011111100110110110: color_data = 12'b111100001111;
20'b00011111100110110111: color_data = 12'b111100001111;
20'b00011111110011100100: color_data = 12'b000000001111;
20'b00011111110011100101: color_data = 12'b000000001111;
20'b00011111110011100110: color_data = 12'b000000001111;
20'b00011111110011100111: color_data = 12'b000000001111;
20'b00011111110011101000: color_data = 12'b000000001111;
20'b00011111110011101001: color_data = 12'b000000001111;
20'b00011111110011101010: color_data = 12'b000000001111;
20'b00011111110011101011: color_data = 12'b000000001111;
20'b00011111110100000101: color_data = 12'b000001101111;
20'b00011111110100000110: color_data = 12'b000001101111;
20'b00011111110100000111: color_data = 12'b000001101111;
20'b00011111110100001000: color_data = 12'b000001101111;
20'b00011111110100001001: color_data = 12'b000001101111;
20'b00011111110100001010: color_data = 12'b000001101111;
20'b00011111110100001011: color_data = 12'b000001101111;
20'b00011111110100001100: color_data = 12'b000001101111;
20'b00011111110100111110: color_data = 12'b000011111111;
20'b00011111110100111111: color_data = 12'b000011111111;
20'b00011111110101000000: color_data = 12'b000011111111;
20'b00011111110101000001: color_data = 12'b000011111111;
20'b00011111110101000010: color_data = 12'b000011111111;
20'b00011111110101000011: color_data = 12'b000011111111;
20'b00011111110101000100: color_data = 12'b000011111111;
20'b00011111110101000101: color_data = 12'b000011111111;
20'b00011111110101011111: color_data = 12'b111101110000;
20'b00011111110101100000: color_data = 12'b111101110000;
20'b00011111110101100001: color_data = 12'b111101110000;
20'b00011111110101100010: color_data = 12'b111101110000;
20'b00011111110101100011: color_data = 12'b111101110000;
20'b00011111110101100100: color_data = 12'b111101110000;
20'b00011111110101100101: color_data = 12'b111101110000;
20'b00011111110101100110: color_data = 12'b111101110000;
20'b00011111110101110111: color_data = 12'b111101100000;
20'b00011111110101111000: color_data = 12'b111101100000;
20'b00011111110101111001: color_data = 12'b111101100000;
20'b00011111110101111010: color_data = 12'b111101100000;
20'b00011111110101111011: color_data = 12'b111101100000;
20'b00011111110101111100: color_data = 12'b111101100000;
20'b00011111110101111101: color_data = 12'b111101100000;
20'b00011111110101111110: color_data = 12'b111101100000;
20'b00011111110110000111: color_data = 12'b000011110000;
20'b00011111110110001000: color_data = 12'b000011110000;
20'b00011111110110001001: color_data = 12'b000011110000;
20'b00011111110110001010: color_data = 12'b000011110000;
20'b00011111110110001011: color_data = 12'b000011110000;
20'b00011111110110001100: color_data = 12'b000011110000;
20'b00011111110110001101: color_data = 12'b000011110000;
20'b00011111110110001110: color_data = 12'b000011110000;
20'b00011111110110001111: color_data = 12'b000011110000;
20'b00011111110110110000: color_data = 12'b111100001111;
20'b00011111110110110001: color_data = 12'b111100001111;
20'b00011111110110110010: color_data = 12'b111100001111;
20'b00011111110110110011: color_data = 12'b111100001111;
20'b00011111110110110100: color_data = 12'b111100001111;
20'b00011111110110110101: color_data = 12'b111100001111;
20'b00011111110110110110: color_data = 12'b111100001111;
20'b00011111110110110111: color_data = 12'b111100001111;
20'b00100000000011100100: color_data = 12'b000000001111;
20'b00100000000011100101: color_data = 12'b000000001111;
20'b00100000000011100110: color_data = 12'b000000001111;
20'b00100000000011100111: color_data = 12'b000000001111;
20'b00100000000011101000: color_data = 12'b000000001111;
20'b00100000000011101001: color_data = 12'b000000001111;
20'b00100000000011101010: color_data = 12'b000000001111;
20'b00100000000011101011: color_data = 12'b000000001111;
20'b00100000000100000101: color_data = 12'b000001101111;
20'b00100000000100000110: color_data = 12'b000001101111;
20'b00100000000100000111: color_data = 12'b000001101111;
20'b00100000000100001000: color_data = 12'b000001101111;
20'b00100000000100001001: color_data = 12'b000001101111;
20'b00100000000100001010: color_data = 12'b000001101111;
20'b00100000000100001011: color_data = 12'b000001101111;
20'b00100000000100001100: color_data = 12'b000001101111;
20'b00100000000100001101: color_data = 12'b000001101111;
20'b00100000000100001110: color_data = 12'b000001101111;
20'b00100000000100001111: color_data = 12'b000001101111;
20'b00100000000100010000: color_data = 12'b000001101111;
20'b00100000000100010001: color_data = 12'b000001101111;
20'b00100000000100010010: color_data = 12'b000001101111;
20'b00100000000100010011: color_data = 12'b000001101111;
20'b00100000000100010100: color_data = 12'b000001101111;
20'b00100000000100010101: color_data = 12'b000001101111;
20'b00100000000100010110: color_data = 12'b000001101111;
20'b00100000000100010111: color_data = 12'b000001101111;
20'b00100000000100011000: color_data = 12'b000001101111;
20'b00100000000100011001: color_data = 12'b000001101111;
20'b00100000000100011010: color_data = 12'b000001101111;
20'b00100000000100011011: color_data = 12'b000001101111;
20'b00100000000100011100: color_data = 12'b000001101111;
20'b00100000000100011101: color_data = 12'b000001101111;
20'b00100000000100011110: color_data = 12'b000001101111;
20'b00100000000100011111: color_data = 12'b000001101111;
20'b00100000000100100000: color_data = 12'b000001101111;
20'b00100000000100100001: color_data = 12'b000001101111;
20'b00100000000100100010: color_data = 12'b000001101111;
20'b00100000000100100011: color_data = 12'b000001101111;
20'b00100000000100100100: color_data = 12'b000001101111;
20'b00100000000100111110: color_data = 12'b000011111111;
20'b00100000000100111111: color_data = 12'b000011111111;
20'b00100000000101000000: color_data = 12'b000011111111;
20'b00100000000101000001: color_data = 12'b000011111111;
20'b00100000000101000010: color_data = 12'b000011111111;
20'b00100000000101000011: color_data = 12'b000011111111;
20'b00100000000101000100: color_data = 12'b000011111111;
20'b00100000000101000101: color_data = 12'b000011111111;
20'b00100000000101011111: color_data = 12'b111101110000;
20'b00100000000101100000: color_data = 12'b111101110000;
20'b00100000000101100001: color_data = 12'b111101110000;
20'b00100000000101100010: color_data = 12'b111101110000;
20'b00100000000101100011: color_data = 12'b111101110000;
20'b00100000000101100100: color_data = 12'b111101110000;
20'b00100000000101100101: color_data = 12'b111101110000;
20'b00100000000101100110: color_data = 12'b111101110000;
20'b00100000000101110111: color_data = 12'b111101100000;
20'b00100000000101111000: color_data = 12'b111101100000;
20'b00100000000101111001: color_data = 12'b111101100000;
20'b00100000000101111010: color_data = 12'b111101100000;
20'b00100000000101111011: color_data = 12'b111101100000;
20'b00100000000101111100: color_data = 12'b111101100000;
20'b00100000000101111101: color_data = 12'b111101100000;
20'b00100000000101111110: color_data = 12'b111101100000;
20'b00100000000110000111: color_data = 12'b000011110000;
20'b00100000000110001000: color_data = 12'b000011110000;
20'b00100000000110001001: color_data = 12'b000011110000;
20'b00100000000110001010: color_data = 12'b000011110000;
20'b00100000000110001011: color_data = 12'b000011110000;
20'b00100000000110001100: color_data = 12'b000011110000;
20'b00100000000110001101: color_data = 12'b000011110000;
20'b00100000000110001110: color_data = 12'b000011110000;
20'b00100000000110001111: color_data = 12'b000011110000;
20'b00100000000110011000: color_data = 12'b111100001111;
20'b00100000000110011001: color_data = 12'b111100001111;
20'b00100000000110011010: color_data = 12'b111100001111;
20'b00100000000110011011: color_data = 12'b111100001111;
20'b00100000000110011100: color_data = 12'b111100001111;
20'b00100000000110011101: color_data = 12'b111100001111;
20'b00100000000110011110: color_data = 12'b111100001111;
20'b00100000000110011111: color_data = 12'b111100001111;
20'b00100000000110100000: color_data = 12'b111100001111;
20'b00100000000110100001: color_data = 12'b111100001111;
20'b00100000000110100010: color_data = 12'b111100001111;
20'b00100000000110100011: color_data = 12'b111100001111;
20'b00100000000110100100: color_data = 12'b111100001111;
20'b00100000000110100101: color_data = 12'b111100001111;
20'b00100000000110100110: color_data = 12'b111100001111;
20'b00100000000110100111: color_data = 12'b111100001111;
20'b00100000000110101000: color_data = 12'b111100001111;
20'b00100000000110101001: color_data = 12'b111100001111;
20'b00100000000110101010: color_data = 12'b111100001111;
20'b00100000000110101011: color_data = 12'b111100001111;
20'b00100000000110101100: color_data = 12'b111100001111;
20'b00100000000110101101: color_data = 12'b111100001111;
20'b00100000000110101110: color_data = 12'b111100001111;
20'b00100000000110101111: color_data = 12'b111100001111;
20'b00100000000110110000: color_data = 12'b111100001111;
20'b00100000000110110001: color_data = 12'b111100001111;
20'b00100000000110110010: color_data = 12'b111100001111;
20'b00100000000110110011: color_data = 12'b111100001111;
20'b00100000000110110100: color_data = 12'b111100001111;
20'b00100000000110110101: color_data = 12'b111100001111;
20'b00100000000110110110: color_data = 12'b111100001111;
20'b00100000000110110111: color_data = 12'b111100001111;
20'b00100000010011100100: color_data = 12'b000000001111;
20'b00100000010011100101: color_data = 12'b000000001111;
20'b00100000010011100110: color_data = 12'b000000001111;
20'b00100000010011100111: color_data = 12'b000000001111;
20'b00100000010011101000: color_data = 12'b000000001111;
20'b00100000010011101001: color_data = 12'b000000001111;
20'b00100000010011101010: color_data = 12'b000000001111;
20'b00100000010011101011: color_data = 12'b000000001111;
20'b00100000010100000101: color_data = 12'b000001101111;
20'b00100000010100000110: color_data = 12'b000001101111;
20'b00100000010100000111: color_data = 12'b000001101111;
20'b00100000010100001000: color_data = 12'b000001101111;
20'b00100000010100001001: color_data = 12'b000001101111;
20'b00100000010100001010: color_data = 12'b000001101111;
20'b00100000010100001011: color_data = 12'b000001101111;
20'b00100000010100001100: color_data = 12'b000001101111;
20'b00100000010100001101: color_data = 12'b000001101111;
20'b00100000010100001110: color_data = 12'b000001101111;
20'b00100000010100001111: color_data = 12'b000001101111;
20'b00100000010100010000: color_data = 12'b000001101111;
20'b00100000010100010001: color_data = 12'b000001101111;
20'b00100000010100010010: color_data = 12'b000001101111;
20'b00100000010100010011: color_data = 12'b000001101111;
20'b00100000010100010100: color_data = 12'b000001101111;
20'b00100000010100010101: color_data = 12'b000001101111;
20'b00100000010100010110: color_data = 12'b000001101111;
20'b00100000010100010111: color_data = 12'b000001101111;
20'b00100000010100011000: color_data = 12'b000001101111;
20'b00100000010100011001: color_data = 12'b000001101111;
20'b00100000010100011010: color_data = 12'b000001101111;
20'b00100000010100011011: color_data = 12'b000001101111;
20'b00100000010100011100: color_data = 12'b000001101111;
20'b00100000010100011101: color_data = 12'b000001101111;
20'b00100000010100011110: color_data = 12'b000001101111;
20'b00100000010100011111: color_data = 12'b000001101111;
20'b00100000010100100000: color_data = 12'b000001101111;
20'b00100000010100100001: color_data = 12'b000001101111;
20'b00100000010100100010: color_data = 12'b000001101111;
20'b00100000010100100011: color_data = 12'b000001101111;
20'b00100000010100100100: color_data = 12'b000001101111;
20'b00100000010100111110: color_data = 12'b000011111111;
20'b00100000010100111111: color_data = 12'b000011111111;
20'b00100000010101000000: color_data = 12'b000011111111;
20'b00100000010101000001: color_data = 12'b000011111111;
20'b00100000010101000010: color_data = 12'b000011111111;
20'b00100000010101000011: color_data = 12'b000011111111;
20'b00100000010101000100: color_data = 12'b000011111111;
20'b00100000010101000101: color_data = 12'b000011111111;
20'b00100000010101011111: color_data = 12'b111101110000;
20'b00100000010101100000: color_data = 12'b111101110000;
20'b00100000010101100001: color_data = 12'b111101110000;
20'b00100000010101100010: color_data = 12'b111101110000;
20'b00100000010101100011: color_data = 12'b111101110000;
20'b00100000010101100100: color_data = 12'b111101110000;
20'b00100000010101100101: color_data = 12'b111101110000;
20'b00100000010101100110: color_data = 12'b111101110000;
20'b00100000010101110111: color_data = 12'b111101100000;
20'b00100000010101111000: color_data = 12'b111101100000;
20'b00100000010101111001: color_data = 12'b111101100000;
20'b00100000010101111010: color_data = 12'b111101100000;
20'b00100000010101111011: color_data = 12'b111101100000;
20'b00100000010101111100: color_data = 12'b111101100000;
20'b00100000010101111101: color_data = 12'b111101100000;
20'b00100000010101111110: color_data = 12'b111101100000;
20'b00100000010110000111: color_data = 12'b000011110000;
20'b00100000010110001000: color_data = 12'b000011110000;
20'b00100000010110001001: color_data = 12'b000011110000;
20'b00100000010110001010: color_data = 12'b000011110000;
20'b00100000010110001011: color_data = 12'b000011110000;
20'b00100000010110001100: color_data = 12'b000011110000;
20'b00100000010110001101: color_data = 12'b000011110000;
20'b00100000010110001110: color_data = 12'b000011110000;
20'b00100000010110001111: color_data = 12'b000011110000;
20'b00100000010110011000: color_data = 12'b111100001111;
20'b00100000010110011001: color_data = 12'b111100001111;
20'b00100000010110011010: color_data = 12'b111100001111;
20'b00100000010110011011: color_data = 12'b111100001111;
20'b00100000010110011100: color_data = 12'b111100001111;
20'b00100000010110011101: color_data = 12'b111100001111;
20'b00100000010110011110: color_data = 12'b111100001111;
20'b00100000010110011111: color_data = 12'b111100001111;
20'b00100000010110100000: color_data = 12'b111100001111;
20'b00100000010110100001: color_data = 12'b111100001111;
20'b00100000010110100010: color_data = 12'b111100001111;
20'b00100000010110100011: color_data = 12'b111100001111;
20'b00100000010110100100: color_data = 12'b111100001111;
20'b00100000010110100101: color_data = 12'b111100001111;
20'b00100000010110100110: color_data = 12'b111100001111;
20'b00100000010110100111: color_data = 12'b111100001111;
20'b00100000010110101000: color_data = 12'b111100001111;
20'b00100000010110101001: color_data = 12'b111100001111;
20'b00100000010110101010: color_data = 12'b111100001111;
20'b00100000010110101011: color_data = 12'b111100001111;
20'b00100000010110101100: color_data = 12'b111100001111;
20'b00100000010110101101: color_data = 12'b111100001111;
20'b00100000010110101110: color_data = 12'b111100001111;
20'b00100000010110101111: color_data = 12'b111100001111;
20'b00100000010110110000: color_data = 12'b111100001111;
20'b00100000010110110001: color_data = 12'b111100001111;
20'b00100000010110110010: color_data = 12'b111100001111;
20'b00100000010110110011: color_data = 12'b111100001111;
20'b00100000010110110100: color_data = 12'b111100001111;
20'b00100000010110110101: color_data = 12'b111100001111;
20'b00100000010110110110: color_data = 12'b111100001111;
20'b00100000010110110111: color_data = 12'b111100001111;
20'b00100000100011100100: color_data = 12'b000000001111;
20'b00100000100011100101: color_data = 12'b000000001111;
20'b00100000100011100110: color_data = 12'b000000001111;
20'b00100000100011100111: color_data = 12'b000000001111;
20'b00100000100011101000: color_data = 12'b000000001111;
20'b00100000100011101001: color_data = 12'b000000001111;
20'b00100000100011101010: color_data = 12'b000000001111;
20'b00100000100011101011: color_data = 12'b000000001111;
20'b00100000100100000101: color_data = 12'b000001101111;
20'b00100000100100000110: color_data = 12'b000001101111;
20'b00100000100100000111: color_data = 12'b000001101111;
20'b00100000100100001000: color_data = 12'b000001101111;
20'b00100000100100001001: color_data = 12'b000001101111;
20'b00100000100100001010: color_data = 12'b000001101111;
20'b00100000100100001011: color_data = 12'b000001101111;
20'b00100000100100001100: color_data = 12'b000001101111;
20'b00100000100100001101: color_data = 12'b000001101111;
20'b00100000100100001110: color_data = 12'b000001101111;
20'b00100000100100001111: color_data = 12'b000001101111;
20'b00100000100100010000: color_data = 12'b000001101111;
20'b00100000100100010001: color_data = 12'b000001101111;
20'b00100000100100010010: color_data = 12'b000001101111;
20'b00100000100100010011: color_data = 12'b000001101111;
20'b00100000100100010100: color_data = 12'b000001101111;
20'b00100000100100010101: color_data = 12'b000001101111;
20'b00100000100100010110: color_data = 12'b000001101111;
20'b00100000100100010111: color_data = 12'b000001101111;
20'b00100000100100011000: color_data = 12'b000001101111;
20'b00100000100100011001: color_data = 12'b000001101111;
20'b00100000100100011010: color_data = 12'b000001101111;
20'b00100000100100011011: color_data = 12'b000001101111;
20'b00100000100100011100: color_data = 12'b000001101111;
20'b00100000100100011101: color_data = 12'b000001101111;
20'b00100000100100011110: color_data = 12'b000001101111;
20'b00100000100100011111: color_data = 12'b000001101111;
20'b00100000100100100000: color_data = 12'b000001101111;
20'b00100000100100100001: color_data = 12'b000001101111;
20'b00100000100100100010: color_data = 12'b000001101111;
20'b00100000100100100011: color_data = 12'b000001101111;
20'b00100000100100100100: color_data = 12'b000001101111;
20'b00100000100100111110: color_data = 12'b000011111111;
20'b00100000100100111111: color_data = 12'b000011111111;
20'b00100000100101000000: color_data = 12'b000011111111;
20'b00100000100101000001: color_data = 12'b000011111111;
20'b00100000100101000010: color_data = 12'b000011111111;
20'b00100000100101000011: color_data = 12'b000011111111;
20'b00100000100101000100: color_data = 12'b000011111111;
20'b00100000100101000101: color_data = 12'b000011111111;
20'b00100000100101011111: color_data = 12'b111101110000;
20'b00100000100101100000: color_data = 12'b111101110000;
20'b00100000100101100001: color_data = 12'b111101110000;
20'b00100000100101100010: color_data = 12'b111101110000;
20'b00100000100101100011: color_data = 12'b111101110000;
20'b00100000100101100100: color_data = 12'b111101110000;
20'b00100000100101100101: color_data = 12'b111101110000;
20'b00100000100101100110: color_data = 12'b111101110000;
20'b00100000100101110111: color_data = 12'b111101100000;
20'b00100000100101111000: color_data = 12'b111101100000;
20'b00100000100101111001: color_data = 12'b111101100000;
20'b00100000100101111010: color_data = 12'b111101100000;
20'b00100000100101111011: color_data = 12'b111101100000;
20'b00100000100101111100: color_data = 12'b111101100000;
20'b00100000100101111101: color_data = 12'b111101100000;
20'b00100000100101111110: color_data = 12'b111101100000;
20'b00100000100110000111: color_data = 12'b000011110000;
20'b00100000100110001000: color_data = 12'b000011110000;
20'b00100000100110001001: color_data = 12'b000011110000;
20'b00100000100110001010: color_data = 12'b000011110000;
20'b00100000100110001011: color_data = 12'b000011110000;
20'b00100000100110001100: color_data = 12'b000011110000;
20'b00100000100110001101: color_data = 12'b000011110000;
20'b00100000100110001110: color_data = 12'b000011110000;
20'b00100000100110001111: color_data = 12'b000011110000;
20'b00100000100110011000: color_data = 12'b111100001111;
20'b00100000100110011001: color_data = 12'b111100001111;
20'b00100000100110011010: color_data = 12'b111100001111;
20'b00100000100110011011: color_data = 12'b111100001111;
20'b00100000100110011100: color_data = 12'b111100001111;
20'b00100000100110011101: color_data = 12'b111100001111;
20'b00100000100110011110: color_data = 12'b111100001111;
20'b00100000100110011111: color_data = 12'b111100001111;
20'b00100000100110100000: color_data = 12'b111100001111;
20'b00100000100110100001: color_data = 12'b111100001111;
20'b00100000100110100010: color_data = 12'b111100001111;
20'b00100000100110100011: color_data = 12'b111100001111;
20'b00100000100110100100: color_data = 12'b111100001111;
20'b00100000100110100101: color_data = 12'b111100001111;
20'b00100000100110100110: color_data = 12'b111100001111;
20'b00100000100110100111: color_data = 12'b111100001111;
20'b00100000100110101000: color_data = 12'b111100001111;
20'b00100000100110101001: color_data = 12'b111100001111;
20'b00100000100110101010: color_data = 12'b111100001111;
20'b00100000100110101011: color_data = 12'b111100001111;
20'b00100000100110101100: color_data = 12'b111100001111;
20'b00100000100110101101: color_data = 12'b111100001111;
20'b00100000100110101110: color_data = 12'b111100001111;
20'b00100000100110101111: color_data = 12'b111100001111;
20'b00100000100110110000: color_data = 12'b111100001111;
20'b00100000100110110001: color_data = 12'b111100001111;
20'b00100000100110110010: color_data = 12'b111100001111;
20'b00100000100110110011: color_data = 12'b111100001111;
20'b00100000100110110100: color_data = 12'b111100001111;
20'b00100000100110110101: color_data = 12'b111100001111;
20'b00100000100110110110: color_data = 12'b111100001111;
20'b00100000100110110111: color_data = 12'b111100001111;
20'b00100000110011100100: color_data = 12'b000000001111;
20'b00100000110011100101: color_data = 12'b000000001111;
20'b00100000110011100110: color_data = 12'b000000001111;
20'b00100000110011100111: color_data = 12'b000000001111;
20'b00100000110011101000: color_data = 12'b000000001111;
20'b00100000110011101001: color_data = 12'b000000001111;
20'b00100000110011101010: color_data = 12'b000000001111;
20'b00100000110011101011: color_data = 12'b000000001111;
20'b00100000110100000101: color_data = 12'b000001101111;
20'b00100000110100000110: color_data = 12'b000001101111;
20'b00100000110100000111: color_data = 12'b000001101111;
20'b00100000110100001000: color_data = 12'b000001101111;
20'b00100000110100001001: color_data = 12'b000001101111;
20'b00100000110100001010: color_data = 12'b000001101111;
20'b00100000110100001011: color_data = 12'b000001101111;
20'b00100000110100001100: color_data = 12'b000001101111;
20'b00100000110100001101: color_data = 12'b000001101111;
20'b00100000110100001110: color_data = 12'b000001101111;
20'b00100000110100001111: color_data = 12'b000001101111;
20'b00100000110100010000: color_data = 12'b000001101111;
20'b00100000110100010001: color_data = 12'b000001101111;
20'b00100000110100010010: color_data = 12'b000001101111;
20'b00100000110100010011: color_data = 12'b000001101111;
20'b00100000110100010100: color_data = 12'b000001101111;
20'b00100000110100010101: color_data = 12'b000001101111;
20'b00100000110100010110: color_data = 12'b000001101111;
20'b00100000110100010111: color_data = 12'b000001101111;
20'b00100000110100011000: color_data = 12'b000001101111;
20'b00100000110100011001: color_data = 12'b000001101111;
20'b00100000110100011010: color_data = 12'b000001101111;
20'b00100000110100011011: color_data = 12'b000001101111;
20'b00100000110100011100: color_data = 12'b000001101111;
20'b00100000110100011101: color_data = 12'b000001101111;
20'b00100000110100011110: color_data = 12'b000001101111;
20'b00100000110100011111: color_data = 12'b000001101111;
20'b00100000110100100000: color_data = 12'b000001101111;
20'b00100000110100100001: color_data = 12'b000001101111;
20'b00100000110100100010: color_data = 12'b000001101111;
20'b00100000110100100011: color_data = 12'b000001101111;
20'b00100000110100100100: color_data = 12'b000001101111;
20'b00100000110100111110: color_data = 12'b000011111111;
20'b00100000110100111111: color_data = 12'b000011111111;
20'b00100000110101000000: color_data = 12'b000011111111;
20'b00100000110101000001: color_data = 12'b000011111111;
20'b00100000110101000010: color_data = 12'b000011111111;
20'b00100000110101000011: color_data = 12'b000011111111;
20'b00100000110101000100: color_data = 12'b000011111111;
20'b00100000110101000101: color_data = 12'b000011111111;
20'b00100000110101011111: color_data = 12'b111101110000;
20'b00100000110101100000: color_data = 12'b111101110000;
20'b00100000110101100001: color_data = 12'b111101110000;
20'b00100000110101100010: color_data = 12'b111101110000;
20'b00100000110101100011: color_data = 12'b111101110000;
20'b00100000110101100100: color_data = 12'b111101110000;
20'b00100000110101100101: color_data = 12'b111101110000;
20'b00100000110101100110: color_data = 12'b111101110000;
20'b00100000110101110111: color_data = 12'b111101100000;
20'b00100000110101111000: color_data = 12'b111101100000;
20'b00100000110101111001: color_data = 12'b111101100000;
20'b00100000110101111010: color_data = 12'b111101100000;
20'b00100000110101111011: color_data = 12'b111101100000;
20'b00100000110101111100: color_data = 12'b111101100000;
20'b00100000110101111101: color_data = 12'b111101100000;
20'b00100000110101111110: color_data = 12'b111101100000;
20'b00100000110110000111: color_data = 12'b000011110000;
20'b00100000110110001000: color_data = 12'b000011110000;
20'b00100000110110001001: color_data = 12'b000011110000;
20'b00100000110110001010: color_data = 12'b000011110000;
20'b00100000110110001011: color_data = 12'b000011110000;
20'b00100000110110001100: color_data = 12'b000011110000;
20'b00100000110110001101: color_data = 12'b000011110000;
20'b00100000110110001110: color_data = 12'b000011110000;
20'b00100000110110001111: color_data = 12'b000011110000;
20'b00100000110110011000: color_data = 12'b111100001111;
20'b00100000110110011001: color_data = 12'b111100001111;
20'b00100000110110011010: color_data = 12'b111100001111;
20'b00100000110110011011: color_data = 12'b111100001111;
20'b00100000110110011100: color_data = 12'b111100001111;
20'b00100000110110011101: color_data = 12'b111100001111;
20'b00100000110110011110: color_data = 12'b111100001111;
20'b00100000110110011111: color_data = 12'b111100001111;
20'b00100000110110100000: color_data = 12'b111100001111;
20'b00100000110110100001: color_data = 12'b111100001111;
20'b00100000110110100010: color_data = 12'b111100001111;
20'b00100000110110100011: color_data = 12'b111100001111;
20'b00100000110110100100: color_data = 12'b111100001111;
20'b00100000110110100101: color_data = 12'b111100001111;
20'b00100000110110100110: color_data = 12'b111100001111;
20'b00100000110110100111: color_data = 12'b111100001111;
20'b00100000110110101000: color_data = 12'b111100001111;
20'b00100000110110101001: color_data = 12'b111100001111;
20'b00100000110110101010: color_data = 12'b111100001111;
20'b00100000110110101011: color_data = 12'b111100001111;
20'b00100000110110101100: color_data = 12'b111100001111;
20'b00100000110110101101: color_data = 12'b111100001111;
20'b00100000110110101110: color_data = 12'b111100001111;
20'b00100000110110101111: color_data = 12'b111100001111;
20'b00100000110110110000: color_data = 12'b111100001111;
20'b00100000110110110001: color_data = 12'b111100001111;
20'b00100000110110110010: color_data = 12'b111100001111;
20'b00100000110110110011: color_data = 12'b111100001111;
20'b00100000110110110100: color_data = 12'b111100001111;
20'b00100000110110110101: color_data = 12'b111100001111;
20'b00100000110110110110: color_data = 12'b111100001111;
20'b00100000110110110111: color_data = 12'b111100001111;
20'b00100001000011100100: color_data = 12'b000000001111;
20'b00100001000011100101: color_data = 12'b000000001111;
20'b00100001000011100110: color_data = 12'b000000001111;
20'b00100001000011100111: color_data = 12'b000000001111;
20'b00100001000011101000: color_data = 12'b000000001111;
20'b00100001000011101001: color_data = 12'b000000001111;
20'b00100001000011101010: color_data = 12'b000000001111;
20'b00100001000011101011: color_data = 12'b000000001111;
20'b00100001000100000101: color_data = 12'b000001101111;
20'b00100001000100000110: color_data = 12'b000001101111;
20'b00100001000100000111: color_data = 12'b000001101111;
20'b00100001000100001000: color_data = 12'b000001101111;
20'b00100001000100001001: color_data = 12'b000001101111;
20'b00100001000100001010: color_data = 12'b000001101111;
20'b00100001000100001011: color_data = 12'b000001101111;
20'b00100001000100001100: color_data = 12'b000001101111;
20'b00100001000100001101: color_data = 12'b000001101111;
20'b00100001000100001110: color_data = 12'b000001101111;
20'b00100001000100001111: color_data = 12'b000001101111;
20'b00100001000100010000: color_data = 12'b000001101111;
20'b00100001000100010001: color_data = 12'b000001101111;
20'b00100001000100010010: color_data = 12'b000001101111;
20'b00100001000100010011: color_data = 12'b000001101111;
20'b00100001000100010100: color_data = 12'b000001101111;
20'b00100001000100010101: color_data = 12'b000001101111;
20'b00100001000100010110: color_data = 12'b000001101111;
20'b00100001000100010111: color_data = 12'b000001101111;
20'b00100001000100011000: color_data = 12'b000001101111;
20'b00100001000100011001: color_data = 12'b000001101111;
20'b00100001000100011010: color_data = 12'b000001101111;
20'b00100001000100011011: color_data = 12'b000001101111;
20'b00100001000100011100: color_data = 12'b000001101111;
20'b00100001000100011101: color_data = 12'b000001101111;
20'b00100001000100011110: color_data = 12'b000001101111;
20'b00100001000100011111: color_data = 12'b000001101111;
20'b00100001000100100000: color_data = 12'b000001101111;
20'b00100001000100100001: color_data = 12'b000001101111;
20'b00100001000100100010: color_data = 12'b000001101111;
20'b00100001000100100011: color_data = 12'b000001101111;
20'b00100001000100100100: color_data = 12'b000001101111;
20'b00100001000100111110: color_data = 12'b000011111111;
20'b00100001000100111111: color_data = 12'b000011111111;
20'b00100001000101000000: color_data = 12'b000011111111;
20'b00100001000101000001: color_data = 12'b000011111111;
20'b00100001000101000010: color_data = 12'b000011111111;
20'b00100001000101000011: color_data = 12'b000011111111;
20'b00100001000101000100: color_data = 12'b000011111111;
20'b00100001000101000101: color_data = 12'b000011111111;
20'b00100001000101011111: color_data = 12'b111101110000;
20'b00100001000101100000: color_data = 12'b111101110000;
20'b00100001000101100001: color_data = 12'b111101110000;
20'b00100001000101100010: color_data = 12'b111101110000;
20'b00100001000101100011: color_data = 12'b111101110000;
20'b00100001000101100100: color_data = 12'b111101110000;
20'b00100001000101100101: color_data = 12'b111101110000;
20'b00100001000101100110: color_data = 12'b111101110000;
20'b00100001000101110111: color_data = 12'b111101100000;
20'b00100001000101111000: color_data = 12'b111101100000;
20'b00100001000101111001: color_data = 12'b111101100000;
20'b00100001000101111010: color_data = 12'b111101100000;
20'b00100001000101111011: color_data = 12'b111101100000;
20'b00100001000101111100: color_data = 12'b111101100000;
20'b00100001000101111101: color_data = 12'b111101100000;
20'b00100001000101111110: color_data = 12'b111101100000;
20'b00100001000110000111: color_data = 12'b000011110000;
20'b00100001000110001000: color_data = 12'b000011110000;
20'b00100001000110001001: color_data = 12'b000011110000;
20'b00100001000110001010: color_data = 12'b000011110000;
20'b00100001000110001011: color_data = 12'b000011110000;
20'b00100001000110001100: color_data = 12'b000011110000;
20'b00100001000110001101: color_data = 12'b000011110000;
20'b00100001000110001110: color_data = 12'b000011110000;
20'b00100001000110001111: color_data = 12'b000011110000;
20'b00100001000110011000: color_data = 12'b111100001111;
20'b00100001000110011001: color_data = 12'b111100001111;
20'b00100001000110011010: color_data = 12'b111100001111;
20'b00100001000110011011: color_data = 12'b111100001111;
20'b00100001000110011100: color_data = 12'b111100001111;
20'b00100001000110011101: color_data = 12'b111100001111;
20'b00100001000110011110: color_data = 12'b111100001111;
20'b00100001000110011111: color_data = 12'b111100001111;
20'b00100001000110100000: color_data = 12'b111100001111;
20'b00100001000110100001: color_data = 12'b111100001111;
20'b00100001000110100010: color_data = 12'b111100001111;
20'b00100001000110100011: color_data = 12'b111100001111;
20'b00100001000110100100: color_data = 12'b111100001111;
20'b00100001000110100101: color_data = 12'b111100001111;
20'b00100001000110100110: color_data = 12'b111100001111;
20'b00100001000110100111: color_data = 12'b111100001111;
20'b00100001000110101000: color_data = 12'b111100001111;
20'b00100001000110101001: color_data = 12'b111100001111;
20'b00100001000110101010: color_data = 12'b111100001111;
20'b00100001000110101011: color_data = 12'b111100001111;
20'b00100001000110101100: color_data = 12'b111100001111;
20'b00100001000110101101: color_data = 12'b111100001111;
20'b00100001000110101110: color_data = 12'b111100001111;
20'b00100001000110101111: color_data = 12'b111100001111;
20'b00100001000110110000: color_data = 12'b111100001111;
20'b00100001000110110001: color_data = 12'b111100001111;
20'b00100001000110110010: color_data = 12'b111100001111;
20'b00100001000110110011: color_data = 12'b111100001111;
20'b00100001000110110100: color_data = 12'b111100001111;
20'b00100001000110110101: color_data = 12'b111100001111;
20'b00100001000110110110: color_data = 12'b111100001111;
20'b00100001000110110111: color_data = 12'b111100001111;
20'b00100001010011100100: color_data = 12'b000000001111;
20'b00100001010011100101: color_data = 12'b000000001111;
20'b00100001010011100110: color_data = 12'b000000001111;
20'b00100001010011100111: color_data = 12'b000000001111;
20'b00100001010011101000: color_data = 12'b000000001111;
20'b00100001010011101001: color_data = 12'b000000001111;
20'b00100001010011101010: color_data = 12'b000000001111;
20'b00100001010011101011: color_data = 12'b000000001111;
20'b00100001010100000101: color_data = 12'b000001101111;
20'b00100001010100000110: color_data = 12'b000001101111;
20'b00100001010100000111: color_data = 12'b000001101111;
20'b00100001010100001000: color_data = 12'b000001101111;
20'b00100001010100001001: color_data = 12'b000001101111;
20'b00100001010100001010: color_data = 12'b000001101111;
20'b00100001010100001011: color_data = 12'b000001101111;
20'b00100001010100001100: color_data = 12'b000001101111;
20'b00100001010100001101: color_data = 12'b000001101111;
20'b00100001010100001110: color_data = 12'b000001101111;
20'b00100001010100001111: color_data = 12'b000001101111;
20'b00100001010100010000: color_data = 12'b000001101111;
20'b00100001010100010001: color_data = 12'b000001101111;
20'b00100001010100010010: color_data = 12'b000001101111;
20'b00100001010100010011: color_data = 12'b000001101111;
20'b00100001010100010100: color_data = 12'b000001101111;
20'b00100001010100010101: color_data = 12'b000001101111;
20'b00100001010100010110: color_data = 12'b000001101111;
20'b00100001010100010111: color_data = 12'b000001101111;
20'b00100001010100011000: color_data = 12'b000001101111;
20'b00100001010100011001: color_data = 12'b000001101111;
20'b00100001010100011010: color_data = 12'b000001101111;
20'b00100001010100011011: color_data = 12'b000001101111;
20'b00100001010100011100: color_data = 12'b000001101111;
20'b00100001010100011101: color_data = 12'b000001101111;
20'b00100001010100011110: color_data = 12'b000001101111;
20'b00100001010100011111: color_data = 12'b000001101111;
20'b00100001010100100000: color_data = 12'b000001101111;
20'b00100001010100100001: color_data = 12'b000001101111;
20'b00100001010100100010: color_data = 12'b000001101111;
20'b00100001010100100011: color_data = 12'b000001101111;
20'b00100001010100100100: color_data = 12'b000001101111;
20'b00100001010100111110: color_data = 12'b000011111111;
20'b00100001010100111111: color_data = 12'b000011111111;
20'b00100001010101000000: color_data = 12'b000011111111;
20'b00100001010101000001: color_data = 12'b000011111111;
20'b00100001010101000010: color_data = 12'b000011111111;
20'b00100001010101000011: color_data = 12'b000011111111;
20'b00100001010101000100: color_data = 12'b000011111111;
20'b00100001010101000101: color_data = 12'b000011111111;
20'b00100001010101011111: color_data = 12'b111101110000;
20'b00100001010101100000: color_data = 12'b111101110000;
20'b00100001010101100001: color_data = 12'b111101110000;
20'b00100001010101100010: color_data = 12'b111101110000;
20'b00100001010101100011: color_data = 12'b111101110000;
20'b00100001010101100100: color_data = 12'b111101110000;
20'b00100001010101100101: color_data = 12'b111101110000;
20'b00100001010101100110: color_data = 12'b111101110000;
20'b00100001010101110111: color_data = 12'b111101100000;
20'b00100001010101111000: color_data = 12'b111101100000;
20'b00100001010101111001: color_data = 12'b111101100000;
20'b00100001010101111010: color_data = 12'b111101100000;
20'b00100001010101111011: color_data = 12'b111101100000;
20'b00100001010101111100: color_data = 12'b111101100000;
20'b00100001010101111101: color_data = 12'b111101100000;
20'b00100001010101111110: color_data = 12'b111101100000;
20'b00100001010110000111: color_data = 12'b000011110000;
20'b00100001010110001000: color_data = 12'b000011110000;
20'b00100001010110001001: color_data = 12'b000011110000;
20'b00100001010110001010: color_data = 12'b000011110000;
20'b00100001010110001011: color_data = 12'b000011110000;
20'b00100001010110001100: color_data = 12'b000011110000;
20'b00100001010110001101: color_data = 12'b000011110000;
20'b00100001010110001110: color_data = 12'b000011110000;
20'b00100001010110001111: color_data = 12'b000011110000;
20'b00100001010110011000: color_data = 12'b111100001111;
20'b00100001010110011001: color_data = 12'b111100001111;
20'b00100001010110011010: color_data = 12'b111100001111;
20'b00100001010110011011: color_data = 12'b111100001111;
20'b00100001010110011100: color_data = 12'b111100001111;
20'b00100001010110011101: color_data = 12'b111100001111;
20'b00100001010110011110: color_data = 12'b111100001111;
20'b00100001010110011111: color_data = 12'b111100001111;
20'b00100001010110100000: color_data = 12'b111100001111;
20'b00100001010110100001: color_data = 12'b111100001111;
20'b00100001010110100010: color_data = 12'b111100001111;
20'b00100001010110100011: color_data = 12'b111100001111;
20'b00100001010110100100: color_data = 12'b111100001111;
20'b00100001010110100101: color_data = 12'b111100001111;
20'b00100001010110100110: color_data = 12'b111100001111;
20'b00100001010110100111: color_data = 12'b111100001111;
20'b00100001010110101000: color_data = 12'b111100001111;
20'b00100001010110101001: color_data = 12'b111100001111;
20'b00100001010110101010: color_data = 12'b111100001111;
20'b00100001010110101011: color_data = 12'b111100001111;
20'b00100001010110101100: color_data = 12'b111100001111;
20'b00100001010110101101: color_data = 12'b111100001111;
20'b00100001010110101110: color_data = 12'b111100001111;
20'b00100001010110101111: color_data = 12'b111100001111;
20'b00100001010110110000: color_data = 12'b111100001111;
20'b00100001010110110001: color_data = 12'b111100001111;
20'b00100001010110110010: color_data = 12'b111100001111;
20'b00100001010110110011: color_data = 12'b111100001111;
20'b00100001010110110100: color_data = 12'b111100001111;
20'b00100001010110110101: color_data = 12'b111100001111;
20'b00100001010110110110: color_data = 12'b111100001111;
20'b00100001010110110111: color_data = 12'b111100001111;
20'b00100001100011100100: color_data = 12'b000000001111;
20'b00100001100011100101: color_data = 12'b000000001111;
20'b00100001100011100110: color_data = 12'b000000001111;
20'b00100001100011100111: color_data = 12'b000000001111;
20'b00100001100011101000: color_data = 12'b000000001111;
20'b00100001100011101001: color_data = 12'b000000001111;
20'b00100001100011101010: color_data = 12'b000000001111;
20'b00100001100011101011: color_data = 12'b000000001111;
20'b00100001100100000101: color_data = 12'b000001101111;
20'b00100001100100000110: color_data = 12'b000001101111;
20'b00100001100100000111: color_data = 12'b000001101111;
20'b00100001100100001000: color_data = 12'b000001101111;
20'b00100001100100001001: color_data = 12'b000001101111;
20'b00100001100100001010: color_data = 12'b000001101111;
20'b00100001100100001011: color_data = 12'b000001101111;
20'b00100001100100001100: color_data = 12'b000001101111;
20'b00100001100100001101: color_data = 12'b000001101111;
20'b00100001100100001110: color_data = 12'b000001101111;
20'b00100001100100001111: color_data = 12'b000001101111;
20'b00100001100100010000: color_data = 12'b000001101111;
20'b00100001100100010001: color_data = 12'b000001101111;
20'b00100001100100010010: color_data = 12'b000001101111;
20'b00100001100100010011: color_data = 12'b000001101111;
20'b00100001100100010100: color_data = 12'b000001101111;
20'b00100001100100010101: color_data = 12'b000001101111;
20'b00100001100100010110: color_data = 12'b000001101111;
20'b00100001100100010111: color_data = 12'b000001101111;
20'b00100001100100011000: color_data = 12'b000001101111;
20'b00100001100100011001: color_data = 12'b000001101111;
20'b00100001100100011010: color_data = 12'b000001101111;
20'b00100001100100011011: color_data = 12'b000001101111;
20'b00100001100100011100: color_data = 12'b000001101111;
20'b00100001100100011101: color_data = 12'b000001101111;
20'b00100001100100011110: color_data = 12'b000001101111;
20'b00100001100100011111: color_data = 12'b000001101111;
20'b00100001100100100000: color_data = 12'b000001101111;
20'b00100001100100100001: color_data = 12'b000001101111;
20'b00100001100100100010: color_data = 12'b000001101111;
20'b00100001100100100011: color_data = 12'b000001101111;
20'b00100001100100100100: color_data = 12'b000001101111;
20'b00100001100100111110: color_data = 12'b000011111111;
20'b00100001100100111111: color_data = 12'b000011111111;
20'b00100001100101000000: color_data = 12'b000011111111;
20'b00100001100101000001: color_data = 12'b000011111111;
20'b00100001100101000010: color_data = 12'b000011111111;
20'b00100001100101000011: color_data = 12'b000011111111;
20'b00100001100101000100: color_data = 12'b000011111111;
20'b00100001100101000101: color_data = 12'b000011111111;
20'b00100001100101011111: color_data = 12'b111101110000;
20'b00100001100101100000: color_data = 12'b111101110000;
20'b00100001100101100001: color_data = 12'b111101110000;
20'b00100001100101100010: color_data = 12'b111101110000;
20'b00100001100101100011: color_data = 12'b111101110000;
20'b00100001100101100100: color_data = 12'b111101110000;
20'b00100001100101100101: color_data = 12'b111101110000;
20'b00100001100101100110: color_data = 12'b111101110000;
20'b00100001100101110111: color_data = 12'b111101100000;
20'b00100001100101111000: color_data = 12'b111101100000;
20'b00100001100101111001: color_data = 12'b111101100000;
20'b00100001100101111010: color_data = 12'b111101100000;
20'b00100001100101111011: color_data = 12'b111101100000;
20'b00100001100101111100: color_data = 12'b111101100000;
20'b00100001100101111101: color_data = 12'b111101100000;
20'b00100001100101111110: color_data = 12'b111101100000;
20'b00100001100110000111: color_data = 12'b000011110000;
20'b00100001100110001000: color_data = 12'b000011110000;
20'b00100001100110001001: color_data = 12'b000011110000;
20'b00100001100110001010: color_data = 12'b000011110000;
20'b00100001100110001011: color_data = 12'b000011110000;
20'b00100001100110001100: color_data = 12'b000011110000;
20'b00100001100110001101: color_data = 12'b000011110000;
20'b00100001100110001110: color_data = 12'b000011110000;
20'b00100001100110001111: color_data = 12'b000011110000;
20'b00100001100110011000: color_data = 12'b111100001111;
20'b00100001100110011001: color_data = 12'b111100001111;
20'b00100001100110011010: color_data = 12'b111100001111;
20'b00100001100110011011: color_data = 12'b111100001111;
20'b00100001100110011100: color_data = 12'b111100001111;
20'b00100001100110011101: color_data = 12'b111100001111;
20'b00100001100110011110: color_data = 12'b111100001111;
20'b00100001100110011111: color_data = 12'b111100001111;
20'b00100001100110100000: color_data = 12'b111100001111;
20'b00100001100110100001: color_data = 12'b111100001111;
20'b00100001100110100010: color_data = 12'b111100001111;
20'b00100001100110100011: color_data = 12'b111100001111;
20'b00100001100110100100: color_data = 12'b111100001111;
20'b00100001100110100101: color_data = 12'b111100001111;
20'b00100001100110100110: color_data = 12'b111100001111;
20'b00100001100110100111: color_data = 12'b111100001111;
20'b00100001100110101000: color_data = 12'b111100001111;
20'b00100001100110101001: color_data = 12'b111100001111;
20'b00100001100110101010: color_data = 12'b111100001111;
20'b00100001100110101011: color_data = 12'b111100001111;
20'b00100001100110101100: color_data = 12'b111100001111;
20'b00100001100110101101: color_data = 12'b111100001111;
20'b00100001100110101110: color_data = 12'b111100001111;
20'b00100001100110101111: color_data = 12'b111100001111;
20'b00100001100110110000: color_data = 12'b111100001111;
20'b00100001100110110001: color_data = 12'b111100001111;
20'b00100001100110110010: color_data = 12'b111100001111;
20'b00100001100110110011: color_data = 12'b111100001111;
20'b00100001100110110100: color_data = 12'b111100001111;
20'b00100001100110110101: color_data = 12'b111100001111;
20'b00100001100110110110: color_data = 12'b111100001111;
20'b00100001100110110111: color_data = 12'b111100001111;
20'b00100001110011100100: color_data = 12'b000000001111;
20'b00100001110011100101: color_data = 12'b000000001111;
20'b00100001110011100110: color_data = 12'b000000001111;
20'b00100001110011100111: color_data = 12'b000000001111;
20'b00100001110011101000: color_data = 12'b000000001111;
20'b00100001110011101001: color_data = 12'b000000001111;
20'b00100001110011101010: color_data = 12'b000000001111;
20'b00100001110011101011: color_data = 12'b000000001111;
20'b00100001110100000101: color_data = 12'b000001101111;
20'b00100001110100000110: color_data = 12'b000001101111;
20'b00100001110100000111: color_data = 12'b000001101111;
20'b00100001110100001000: color_data = 12'b000001101111;
20'b00100001110100001001: color_data = 12'b000001101111;
20'b00100001110100001010: color_data = 12'b000001101111;
20'b00100001110100001011: color_data = 12'b000001101111;
20'b00100001110100001100: color_data = 12'b000001101111;
20'b00100001110100001101: color_data = 12'b000001101111;
20'b00100001110100001110: color_data = 12'b000001101111;
20'b00100001110100001111: color_data = 12'b000001101111;
20'b00100001110100010000: color_data = 12'b000001101111;
20'b00100001110100010001: color_data = 12'b000001101111;
20'b00100001110100010010: color_data = 12'b000001101111;
20'b00100001110100010011: color_data = 12'b000001101111;
20'b00100001110100010100: color_data = 12'b000001101111;
20'b00100001110100010101: color_data = 12'b000001101111;
20'b00100001110100010110: color_data = 12'b000001101111;
20'b00100001110100010111: color_data = 12'b000001101111;
20'b00100001110100011000: color_data = 12'b000001101111;
20'b00100001110100011001: color_data = 12'b000001101111;
20'b00100001110100011010: color_data = 12'b000001101111;
20'b00100001110100011011: color_data = 12'b000001101111;
20'b00100001110100011100: color_data = 12'b000001101111;
20'b00100001110100011101: color_data = 12'b000001101111;
20'b00100001110100011110: color_data = 12'b000001101111;
20'b00100001110100011111: color_data = 12'b000001101111;
20'b00100001110100100000: color_data = 12'b000001101111;
20'b00100001110100100001: color_data = 12'b000001101111;
20'b00100001110100100010: color_data = 12'b000001101111;
20'b00100001110100100011: color_data = 12'b000001101111;
20'b00100001110100100100: color_data = 12'b000001101111;
20'b00100001110100111110: color_data = 12'b000011111111;
20'b00100001110100111111: color_data = 12'b000011111111;
20'b00100001110101000000: color_data = 12'b000011111111;
20'b00100001110101000001: color_data = 12'b000011111111;
20'b00100001110101000010: color_data = 12'b000011111111;
20'b00100001110101000011: color_data = 12'b000011111111;
20'b00100001110101000100: color_data = 12'b000011111111;
20'b00100001110101000101: color_data = 12'b000011111111;
20'b00100001110101011111: color_data = 12'b111101110000;
20'b00100001110101100000: color_data = 12'b111101110000;
20'b00100001110101100001: color_data = 12'b111101110000;
20'b00100001110101100010: color_data = 12'b111101110000;
20'b00100001110101100011: color_data = 12'b111101110000;
20'b00100001110101100100: color_data = 12'b111101110000;
20'b00100001110101100101: color_data = 12'b111101110000;
20'b00100001110101100110: color_data = 12'b111101110000;
20'b00100001110101110111: color_data = 12'b111101100000;
20'b00100001110101111000: color_data = 12'b111101100000;
20'b00100001110101111001: color_data = 12'b111101100000;
20'b00100001110101111010: color_data = 12'b111101100000;
20'b00100001110101111011: color_data = 12'b111101100000;
20'b00100001110101111100: color_data = 12'b111101100000;
20'b00100001110101111101: color_data = 12'b111101100000;
20'b00100001110101111110: color_data = 12'b111101100000;
20'b00100001110110000111: color_data = 12'b000011110000;
20'b00100001110110001000: color_data = 12'b000011110000;
20'b00100001110110001001: color_data = 12'b000011110000;
20'b00100001110110001010: color_data = 12'b000011110000;
20'b00100001110110001011: color_data = 12'b000011110000;
20'b00100001110110001100: color_data = 12'b000011110000;
20'b00100001110110001101: color_data = 12'b000011110000;
20'b00100001110110001110: color_data = 12'b000011110000;
20'b00100001110110001111: color_data = 12'b000011110000;
20'b00100001110110011000: color_data = 12'b111100001111;
20'b00100001110110011001: color_data = 12'b111100001111;
20'b00100001110110011010: color_data = 12'b111100001111;
20'b00100001110110011011: color_data = 12'b111100001111;
20'b00100001110110011100: color_data = 12'b111100001111;
20'b00100001110110011101: color_data = 12'b111100001111;
20'b00100001110110011110: color_data = 12'b111100001111;
20'b00100001110110011111: color_data = 12'b111100001111;
20'b00100001110110100000: color_data = 12'b111100001111;
20'b00100001110110100001: color_data = 12'b111100001111;
20'b00100001110110100010: color_data = 12'b111100001111;
20'b00100001110110100011: color_data = 12'b111100001111;
20'b00100001110110100100: color_data = 12'b111100001111;
20'b00100001110110100101: color_data = 12'b111100001111;
20'b00100001110110100110: color_data = 12'b111100001111;
20'b00100001110110100111: color_data = 12'b111100001111;
20'b00100001110110101000: color_data = 12'b111100001111;
20'b00100001110110101001: color_data = 12'b111100001111;
20'b00100001110110101010: color_data = 12'b111100001111;
20'b00100001110110101011: color_data = 12'b111100001111;
20'b00100001110110101100: color_data = 12'b111100001111;
20'b00100001110110101101: color_data = 12'b111100001111;
20'b00100001110110101110: color_data = 12'b111100001111;
20'b00100001110110101111: color_data = 12'b111100001111;
20'b00100001110110110000: color_data = 12'b111100001111;
20'b00100001110110110001: color_data = 12'b111100001111;
20'b00100001110110110010: color_data = 12'b111100001111;
20'b00100001110110110011: color_data = 12'b111100001111;
20'b00100001110110110100: color_data = 12'b111100001111;
20'b00100001110110110101: color_data = 12'b111100001111;
20'b00100001110110110110: color_data = 12'b111100001111;
20'b00100001110110110111: color_data = 12'b111100001111;
20'b00100010000011100100: color_data = 12'b000000001111;
20'b00100010000011100101: color_data = 12'b000000001111;
20'b00100010000011100110: color_data = 12'b000000001111;
20'b00100010000011100111: color_data = 12'b000000001111;
20'b00100010000011101000: color_data = 12'b000000001111;
20'b00100010000011101001: color_data = 12'b000000001111;
20'b00100010000011101010: color_data = 12'b000000001111;
20'b00100010000011101011: color_data = 12'b000000001111;
20'b00100010000100000101: color_data = 12'b000001101111;
20'b00100010000100000110: color_data = 12'b000001101111;
20'b00100010000100000111: color_data = 12'b000001101111;
20'b00100010000100001000: color_data = 12'b000001101111;
20'b00100010000100001001: color_data = 12'b000001101111;
20'b00100010000100001010: color_data = 12'b000001101111;
20'b00100010000100001011: color_data = 12'b000001101111;
20'b00100010000100001100: color_data = 12'b000001101111;
20'b00100010000100001101: color_data = 12'b000001101111;
20'b00100010000100001110: color_data = 12'b000001101111;
20'b00100010000100001111: color_data = 12'b000001101111;
20'b00100010000100010000: color_data = 12'b000001101111;
20'b00100010000100010001: color_data = 12'b000001101111;
20'b00100010000100010010: color_data = 12'b000001101111;
20'b00100010000100010011: color_data = 12'b000001101111;
20'b00100010000100010100: color_data = 12'b000001101111;
20'b00100010000100010101: color_data = 12'b000001101111;
20'b00100010000100010110: color_data = 12'b000001101111;
20'b00100010000100010111: color_data = 12'b000001101111;
20'b00100010000100011000: color_data = 12'b000001101111;
20'b00100010000100011001: color_data = 12'b000001101111;
20'b00100010000100011010: color_data = 12'b000001101111;
20'b00100010000100011011: color_data = 12'b000001101111;
20'b00100010000100011100: color_data = 12'b000001101111;
20'b00100010000100011101: color_data = 12'b000001101111;
20'b00100010000100011110: color_data = 12'b000001101111;
20'b00100010000100011111: color_data = 12'b000001101111;
20'b00100010000100100000: color_data = 12'b000001101111;
20'b00100010000100100001: color_data = 12'b000001101111;
20'b00100010000100100010: color_data = 12'b000001101111;
20'b00100010000100100011: color_data = 12'b000001101111;
20'b00100010000100100100: color_data = 12'b000001101111;
20'b00100010000100111110: color_data = 12'b000011111111;
20'b00100010000100111111: color_data = 12'b000011111111;
20'b00100010000101000000: color_data = 12'b000011111111;
20'b00100010000101000001: color_data = 12'b000011111111;
20'b00100010000101000010: color_data = 12'b000011111111;
20'b00100010000101000011: color_data = 12'b000011111111;
20'b00100010000101000100: color_data = 12'b000011111111;
20'b00100010000101000101: color_data = 12'b000011111111;
20'b00100010000101011111: color_data = 12'b111101110000;
20'b00100010000101100000: color_data = 12'b111101110000;
20'b00100010000101100001: color_data = 12'b111101110000;
20'b00100010000101100010: color_data = 12'b111101110000;
20'b00100010000101100011: color_data = 12'b111101110000;
20'b00100010000101100100: color_data = 12'b111101110000;
20'b00100010000101100101: color_data = 12'b111101110000;
20'b00100010000101100110: color_data = 12'b111101110000;
20'b00100010000101110111: color_data = 12'b111101100000;
20'b00100010000101111000: color_data = 12'b111101100000;
20'b00100010000101111001: color_data = 12'b111101100000;
20'b00100010000101111010: color_data = 12'b111101100000;
20'b00100010000101111011: color_data = 12'b111101100000;
20'b00100010000101111100: color_data = 12'b111101100000;
20'b00100010000101111101: color_data = 12'b111101100000;
20'b00100010000101111110: color_data = 12'b111101100000;
20'b00100010000110000111: color_data = 12'b000011110000;
20'b00100010000110001000: color_data = 12'b000011110000;
20'b00100010000110001001: color_data = 12'b000011110000;
20'b00100010000110001010: color_data = 12'b000011110000;
20'b00100010000110001011: color_data = 12'b000011110000;
20'b00100010000110001100: color_data = 12'b000011110000;
20'b00100010000110001101: color_data = 12'b000011110000;
20'b00100010000110001110: color_data = 12'b000011110000;
20'b00100010000110001111: color_data = 12'b000011110000;
20'b00100010000110011000: color_data = 12'b111100001111;
20'b00100010000110011001: color_data = 12'b111100001111;
20'b00100010000110011010: color_data = 12'b111100001111;
20'b00100010000110011011: color_data = 12'b111100001111;
20'b00100010000110011100: color_data = 12'b111100001111;
20'b00100010000110011101: color_data = 12'b111100001111;
20'b00100010000110011110: color_data = 12'b111100001111;
20'b00100010000110011111: color_data = 12'b111100001111;
20'b00100010000110100000: color_data = 12'b111100001111;
20'b00100010000110100001: color_data = 12'b111100001111;
20'b00100010000110100010: color_data = 12'b111100001111;
20'b00100010000110100011: color_data = 12'b111100001111;
20'b00100010000110100100: color_data = 12'b111100001111;
20'b00100010000110100101: color_data = 12'b111100001111;
20'b00100010000110100110: color_data = 12'b111100001111;
20'b00100010000110100111: color_data = 12'b111100001111;
20'b00100010000110101000: color_data = 12'b111100001111;
20'b00100010000110101001: color_data = 12'b111100001111;
20'b00100010000110101010: color_data = 12'b111100001111;
20'b00100010000110101011: color_data = 12'b111100001111;
20'b00100010000110101100: color_data = 12'b111100001111;
20'b00100010000110101101: color_data = 12'b111100001111;
20'b00100010000110101110: color_data = 12'b111100001111;
20'b00100010000110101111: color_data = 12'b111100001111;
20'b00100010000110110000: color_data = 12'b111100001111;
20'b00100010000110110001: color_data = 12'b111100001111;
20'b00100010000110110010: color_data = 12'b111100001111;
20'b00100010000110110011: color_data = 12'b111100001111;
20'b00100010000110110100: color_data = 12'b111100001111;
20'b00100010000110110101: color_data = 12'b111100001111;
20'b00100010000110110110: color_data = 12'b111100001111;
20'b00100010000110110111: color_data = 12'b111100001111;
20'b00100010010011100100: color_data = 12'b000000001111;
20'b00100010010011100101: color_data = 12'b000000001111;
20'b00100010010011100110: color_data = 12'b000000001111;
20'b00100010010011100111: color_data = 12'b000000001111;
20'b00100010010011101000: color_data = 12'b000000001111;
20'b00100010010011101001: color_data = 12'b000000001111;
20'b00100010010011101010: color_data = 12'b000000001111;
20'b00100010010011101011: color_data = 12'b000000001111;
20'b00100010010100000101: color_data = 12'b000001101111;
20'b00100010010100000110: color_data = 12'b000001101111;
20'b00100010010100000111: color_data = 12'b000001101111;
20'b00100010010100001000: color_data = 12'b000001101111;
20'b00100010010100001001: color_data = 12'b000001101111;
20'b00100010010100001010: color_data = 12'b000001101111;
20'b00100010010100001011: color_data = 12'b000001101111;
20'b00100010010100001100: color_data = 12'b000001101111;
20'b00100010010100001101: color_data = 12'b000001101111;
20'b00100010010100001110: color_data = 12'b000001101111;
20'b00100010010100001111: color_data = 12'b000001101111;
20'b00100010010100010000: color_data = 12'b000001101111;
20'b00100010010100010001: color_data = 12'b000001101111;
20'b00100010010100010010: color_data = 12'b000001101111;
20'b00100010010100010011: color_data = 12'b000001101111;
20'b00100010010100010100: color_data = 12'b000001101111;
20'b00100010010100010101: color_data = 12'b000001101111;
20'b00100010010100010110: color_data = 12'b000001101111;
20'b00100010010100010111: color_data = 12'b000001101111;
20'b00100010010100011000: color_data = 12'b000001101111;
20'b00100010010100011001: color_data = 12'b000001101111;
20'b00100010010100011010: color_data = 12'b000001101111;
20'b00100010010100011011: color_data = 12'b000001101111;
20'b00100010010100011100: color_data = 12'b000001101111;
20'b00100010010100011101: color_data = 12'b000001101111;
20'b00100010010100011110: color_data = 12'b000001101111;
20'b00100010010100011111: color_data = 12'b000001101111;
20'b00100010010100100000: color_data = 12'b000001101111;
20'b00100010010100100001: color_data = 12'b000001101111;
20'b00100010010100100010: color_data = 12'b000001101111;
20'b00100010010100100011: color_data = 12'b000001101111;
20'b00100010010100100100: color_data = 12'b000001101111;
20'b00100010010100111110: color_data = 12'b000011111111;
20'b00100010010100111111: color_data = 12'b000011111111;
20'b00100010010101000000: color_data = 12'b000011111111;
20'b00100010010101000001: color_data = 12'b000011111111;
20'b00100010010101000010: color_data = 12'b000011111111;
20'b00100010010101000011: color_data = 12'b000011111111;
20'b00100010010101000100: color_data = 12'b000011111111;
20'b00100010010101000101: color_data = 12'b000011111111;
20'b00100010010101011111: color_data = 12'b111101110000;
20'b00100010010101100000: color_data = 12'b111101110000;
20'b00100010010101100001: color_data = 12'b111101110000;
20'b00100010010101100010: color_data = 12'b111101110000;
20'b00100010010101100011: color_data = 12'b111101110000;
20'b00100010010101100100: color_data = 12'b111101110000;
20'b00100010010101100101: color_data = 12'b111101110000;
20'b00100010010101100110: color_data = 12'b111101110000;
20'b00100010010101110111: color_data = 12'b111101100000;
20'b00100010010101111000: color_data = 12'b111101100000;
20'b00100010010101111001: color_data = 12'b111101100000;
20'b00100010010101111010: color_data = 12'b111101100000;
20'b00100010010101111011: color_data = 12'b111101100000;
20'b00100010010101111100: color_data = 12'b111101100000;
20'b00100010010101111101: color_data = 12'b111101100000;
20'b00100010010101111110: color_data = 12'b111101100000;
20'b00100010010110000111: color_data = 12'b000011110000;
20'b00100010010110001000: color_data = 12'b000011110000;
20'b00100010010110001001: color_data = 12'b000011110000;
20'b00100010010110001010: color_data = 12'b000011110000;
20'b00100010010110001011: color_data = 12'b000011110000;
20'b00100010010110001100: color_data = 12'b000011110000;
20'b00100010010110001101: color_data = 12'b000011110000;
20'b00100010010110001110: color_data = 12'b000011110000;
20'b00100010010110001111: color_data = 12'b000011110000;
20'b00100010010110011000: color_data = 12'b111100001111;
20'b00100010010110011001: color_data = 12'b111100001111;
20'b00100010010110011010: color_data = 12'b111100001111;
20'b00100010010110011011: color_data = 12'b111100001111;
20'b00100010010110011100: color_data = 12'b111100001111;
20'b00100010010110011101: color_data = 12'b111100001111;
20'b00100010010110011110: color_data = 12'b111100001111;
20'b00100010010110011111: color_data = 12'b111100001111;
20'b00100010010110100000: color_data = 12'b111100001111;
20'b00100010010110100001: color_data = 12'b111100001111;
20'b00100010010110100010: color_data = 12'b111100001111;
20'b00100010010110100011: color_data = 12'b111100001111;
20'b00100010010110100100: color_data = 12'b111100001111;
20'b00100010010110100101: color_data = 12'b111100001111;
20'b00100010010110100110: color_data = 12'b111100001111;
20'b00100010010110100111: color_data = 12'b111100001111;
20'b00100010010110101000: color_data = 12'b111100001111;
20'b00100010010110101001: color_data = 12'b111100001111;
20'b00100010010110101010: color_data = 12'b111100001111;
20'b00100010010110101011: color_data = 12'b111100001111;
20'b00100010010110101100: color_data = 12'b111100001111;
20'b00100010010110101101: color_data = 12'b111100001111;
20'b00100010010110101110: color_data = 12'b111100001111;
20'b00100010010110101111: color_data = 12'b111100001111;
20'b00100010010110110000: color_data = 12'b111100001111;
20'b00100010010110110001: color_data = 12'b111100001111;
20'b00100010010110110010: color_data = 12'b111100001111;
20'b00100010010110110011: color_data = 12'b111100001111;
20'b00100010010110110100: color_data = 12'b111100001111;
20'b00100010010110110101: color_data = 12'b111100001111;
20'b00100010010110110110: color_data = 12'b111100001111;
20'b00100010010110110111: color_data = 12'b111100001111;
20'b00100010100011100100: color_data = 12'b000000001111;
20'b00100010100011100101: color_data = 12'b000000001111;
20'b00100010100011100110: color_data = 12'b000000001111;
20'b00100010100011100111: color_data = 12'b000000001111;
20'b00100010100011101000: color_data = 12'b000000001111;
20'b00100010100011101001: color_data = 12'b000000001111;
20'b00100010100011101010: color_data = 12'b000000001111;
20'b00100010100011101011: color_data = 12'b000000001111;
20'b00100010100100000101: color_data = 12'b000001101111;
20'b00100010100100000110: color_data = 12'b000001101111;
20'b00100010100100000111: color_data = 12'b000001101111;
20'b00100010100100001000: color_data = 12'b000001101111;
20'b00100010100100001001: color_data = 12'b000001101111;
20'b00100010100100001010: color_data = 12'b000001101111;
20'b00100010100100001011: color_data = 12'b000001101111;
20'b00100010100100001100: color_data = 12'b000001101111;
20'b00100010100100001101: color_data = 12'b000001101111;
20'b00100010100100001110: color_data = 12'b000001101111;
20'b00100010100100001111: color_data = 12'b000001101111;
20'b00100010100100010000: color_data = 12'b000001101111;
20'b00100010100100010001: color_data = 12'b000001101111;
20'b00100010100100010010: color_data = 12'b000001101111;
20'b00100010100100010011: color_data = 12'b000001101111;
20'b00100010100100010100: color_data = 12'b000001101111;
20'b00100010100100010101: color_data = 12'b000001101111;
20'b00100010100100010110: color_data = 12'b000001101111;
20'b00100010100100010111: color_data = 12'b000001101111;
20'b00100010100100011000: color_data = 12'b000001101111;
20'b00100010100100011001: color_data = 12'b000001101111;
20'b00100010100100011010: color_data = 12'b000001101111;
20'b00100010100100011011: color_data = 12'b000001101111;
20'b00100010100100011100: color_data = 12'b000001101111;
20'b00100010100100011101: color_data = 12'b000001101111;
20'b00100010100100011110: color_data = 12'b000001101111;
20'b00100010100100011111: color_data = 12'b000001101111;
20'b00100010100100100000: color_data = 12'b000001101111;
20'b00100010100100100001: color_data = 12'b000001101111;
20'b00100010100100100010: color_data = 12'b000001101111;
20'b00100010100100100011: color_data = 12'b000001101111;
20'b00100010100100100100: color_data = 12'b000001101111;
20'b00100010100100111110: color_data = 12'b000011111111;
20'b00100010100100111111: color_data = 12'b000011111111;
20'b00100010100101000000: color_data = 12'b000011111111;
20'b00100010100101000001: color_data = 12'b000011111111;
20'b00100010100101000010: color_data = 12'b000011111111;
20'b00100010100101000011: color_data = 12'b000011111111;
20'b00100010100101000100: color_data = 12'b000011111111;
20'b00100010100101000101: color_data = 12'b000011111111;
20'b00100010100101011111: color_data = 12'b111101110000;
20'b00100010100101100000: color_data = 12'b111101110000;
20'b00100010100101100001: color_data = 12'b111101110000;
20'b00100010100101100010: color_data = 12'b111101110000;
20'b00100010100101100011: color_data = 12'b111101110000;
20'b00100010100101100100: color_data = 12'b111101110000;
20'b00100010100101100101: color_data = 12'b111101110000;
20'b00100010100101100110: color_data = 12'b111101110000;
20'b00100010100101110111: color_data = 12'b111101100000;
20'b00100010100101111000: color_data = 12'b111101100000;
20'b00100010100101111001: color_data = 12'b111101100000;
20'b00100010100101111010: color_data = 12'b111101100000;
20'b00100010100101111011: color_data = 12'b111101100000;
20'b00100010100101111100: color_data = 12'b111101100000;
20'b00100010100101111101: color_data = 12'b111101100000;
20'b00100010100101111110: color_data = 12'b111101100000;
20'b00100010100110000111: color_data = 12'b000011110000;
20'b00100010100110001000: color_data = 12'b000011110000;
20'b00100010100110001001: color_data = 12'b000011110000;
20'b00100010100110001010: color_data = 12'b000011110000;
20'b00100010100110001011: color_data = 12'b000011110000;
20'b00100010100110001100: color_data = 12'b000011110000;
20'b00100010100110001101: color_data = 12'b000011110000;
20'b00100010100110001110: color_data = 12'b000011110000;
20'b00100010100110001111: color_data = 12'b000011110000;
20'b00100010100110011000: color_data = 12'b111100001111;
20'b00100010100110011001: color_data = 12'b111100001111;
20'b00100010100110011010: color_data = 12'b111100001111;
20'b00100010100110011011: color_data = 12'b111100001111;
20'b00100010100110011100: color_data = 12'b111100001111;
20'b00100010100110011101: color_data = 12'b111100001111;
20'b00100010100110011110: color_data = 12'b111100001111;
20'b00100010100110011111: color_data = 12'b111100001111;
20'b00100010100110100000: color_data = 12'b111100001111;
20'b00100010100110100001: color_data = 12'b111100001111;
20'b00100010100110100010: color_data = 12'b111100001111;
20'b00100010100110100011: color_data = 12'b111100001111;
20'b00100010100110100100: color_data = 12'b111100001111;
20'b00100010100110100101: color_data = 12'b111100001111;
20'b00100010100110100110: color_data = 12'b111100001111;
20'b00100010100110100111: color_data = 12'b111100001111;
20'b00100010100110101000: color_data = 12'b111100001111;
20'b00100010100110101001: color_data = 12'b111100001111;
20'b00100010100110101010: color_data = 12'b111100001111;
20'b00100010100110101011: color_data = 12'b111100001111;
20'b00100010100110101100: color_data = 12'b111100001111;
20'b00100010100110101101: color_data = 12'b111100001111;
20'b00100010100110101110: color_data = 12'b111100001111;
20'b00100010100110101111: color_data = 12'b111100001111;
20'b00100010100110110000: color_data = 12'b111100001111;
20'b00100010100110110001: color_data = 12'b111100001111;
20'b00100010100110110010: color_data = 12'b111100001111;
20'b00100010100110110011: color_data = 12'b111100001111;
20'b00100010100110110100: color_data = 12'b111100001111;
20'b00100010100110110101: color_data = 12'b111100001111;
20'b00100010100110110110: color_data = 12'b111100001111;
20'b00100010100110110111: color_data = 12'b111100001111;
20'b00100010110011100100: color_data = 12'b000000001111;
20'b00100010110011100101: color_data = 12'b000000001111;
20'b00100010110011100110: color_data = 12'b000000001111;
20'b00100010110011100111: color_data = 12'b000000001111;
20'b00100010110011101000: color_data = 12'b000000001111;
20'b00100010110011101001: color_data = 12'b000000001111;
20'b00100010110011101010: color_data = 12'b000000001111;
20'b00100010110011101011: color_data = 12'b000000001111;
20'b00100010110100000101: color_data = 12'b000001101111;
20'b00100010110100000110: color_data = 12'b000001101111;
20'b00100010110100000111: color_data = 12'b000001101111;
20'b00100010110100001000: color_data = 12'b000001101111;
20'b00100010110100001001: color_data = 12'b000001101111;
20'b00100010110100001010: color_data = 12'b000001101111;
20'b00100010110100001011: color_data = 12'b000001101111;
20'b00100010110100001100: color_data = 12'b000001101111;
20'b00100010110100001101: color_data = 12'b000001101111;
20'b00100010110100001110: color_data = 12'b000001101111;
20'b00100010110100001111: color_data = 12'b000001101111;
20'b00100010110100010000: color_data = 12'b000001101111;
20'b00100010110100010001: color_data = 12'b000001101111;
20'b00100010110100010010: color_data = 12'b000001101111;
20'b00100010110100010011: color_data = 12'b000001101111;
20'b00100010110100010100: color_data = 12'b000001101111;
20'b00100010110100010101: color_data = 12'b000001101111;
20'b00100010110100010110: color_data = 12'b000001101111;
20'b00100010110100010111: color_data = 12'b000001101111;
20'b00100010110100011000: color_data = 12'b000001101111;
20'b00100010110100011001: color_data = 12'b000001101111;
20'b00100010110100011010: color_data = 12'b000001101111;
20'b00100010110100011011: color_data = 12'b000001101111;
20'b00100010110100011100: color_data = 12'b000001101111;
20'b00100010110100011101: color_data = 12'b000001101111;
20'b00100010110100011110: color_data = 12'b000001101111;
20'b00100010110100011111: color_data = 12'b000001101111;
20'b00100010110100100000: color_data = 12'b000001101111;
20'b00100010110100100001: color_data = 12'b000001101111;
20'b00100010110100100010: color_data = 12'b000001101111;
20'b00100010110100100011: color_data = 12'b000001101111;
20'b00100010110100100100: color_data = 12'b000001101111;
20'b00100010110100111110: color_data = 12'b000011111111;
20'b00100010110100111111: color_data = 12'b000011111111;
20'b00100010110101000000: color_data = 12'b000011111111;
20'b00100010110101000001: color_data = 12'b000011111111;
20'b00100010110101000010: color_data = 12'b000011111111;
20'b00100010110101000011: color_data = 12'b000011111111;
20'b00100010110101000100: color_data = 12'b000011111111;
20'b00100010110101000101: color_data = 12'b000011111111;
20'b00100010110101011111: color_data = 12'b111101110000;
20'b00100010110101100000: color_data = 12'b111101110000;
20'b00100010110101100001: color_data = 12'b111101110000;
20'b00100010110101100010: color_data = 12'b111101110000;
20'b00100010110101100011: color_data = 12'b111101110000;
20'b00100010110101100100: color_data = 12'b111101110000;
20'b00100010110101100101: color_data = 12'b111101110000;
20'b00100010110101100110: color_data = 12'b111101110000;
20'b00100010110101110111: color_data = 12'b111101100000;
20'b00100010110101111000: color_data = 12'b111101100000;
20'b00100010110101111001: color_data = 12'b111101100000;
20'b00100010110101111010: color_data = 12'b111101100000;
20'b00100010110101111011: color_data = 12'b111101100000;
20'b00100010110101111100: color_data = 12'b111101100000;
20'b00100010110101111101: color_data = 12'b111101100000;
20'b00100010110101111110: color_data = 12'b111101100000;
20'b00100010110110000111: color_data = 12'b000011110000;
20'b00100010110110001000: color_data = 12'b000011110000;
20'b00100010110110001001: color_data = 12'b000011110000;
20'b00100010110110001010: color_data = 12'b000011110000;
20'b00100010110110001011: color_data = 12'b000011110000;
20'b00100010110110001100: color_data = 12'b000011110000;
20'b00100010110110001101: color_data = 12'b000011110000;
20'b00100010110110001110: color_data = 12'b000011110000;
20'b00100010110110001111: color_data = 12'b000011110000;
20'b00100010110110011000: color_data = 12'b111100001111;
20'b00100010110110011001: color_data = 12'b111100001111;
20'b00100010110110011010: color_data = 12'b111100001111;
20'b00100010110110011011: color_data = 12'b111100001111;
20'b00100010110110011100: color_data = 12'b111100001111;
20'b00100010110110011101: color_data = 12'b111100001111;
20'b00100010110110011110: color_data = 12'b111100001111;
20'b00100010110110011111: color_data = 12'b111100001111;
20'b00100010110110100000: color_data = 12'b111100001111;
20'b00100010110110100001: color_data = 12'b111100001111;
20'b00100010110110100010: color_data = 12'b111100001111;
20'b00100010110110100011: color_data = 12'b111100001111;
20'b00100010110110100100: color_data = 12'b111100001111;
20'b00100010110110100101: color_data = 12'b111100001111;
20'b00100010110110100110: color_data = 12'b111100001111;
20'b00100010110110100111: color_data = 12'b111100001111;
20'b00100010110110101000: color_data = 12'b111100001111;
20'b00100010110110101001: color_data = 12'b111100001111;
20'b00100010110110101010: color_data = 12'b111100001111;
20'b00100010110110101011: color_data = 12'b111100001111;
20'b00100010110110101100: color_data = 12'b111100001111;
20'b00100010110110101101: color_data = 12'b111100001111;
20'b00100010110110101110: color_data = 12'b111100001111;
20'b00100010110110101111: color_data = 12'b111100001111;
20'b00100010110110110000: color_data = 12'b111100001111;
20'b00100010110110110001: color_data = 12'b111100001111;
20'b00100010110110110010: color_data = 12'b111100001111;
20'b00100010110110110011: color_data = 12'b111100001111;
20'b00100010110110110100: color_data = 12'b111100001111;
20'b00100010110110110101: color_data = 12'b111100001111;
20'b00100010110110110110: color_data = 12'b111100001111;
20'b00100010110110110111: color_data = 12'b111100001111;
20'b00110000100100011100: color_data = 12'b111111111111;
20'b00110000100100011101: color_data = 12'b111111111111;
20'b00110000100100011110: color_data = 12'b111111111111;
20'b00110000100100011111: color_data = 12'b111111111111;
20'b00110000100100110000: color_data = 12'b111111111111;
20'b00110000100100110001: color_data = 12'b111111111111;
20'b00110000100100110010: color_data = 12'b111111111111;
20'b00110000100100110011: color_data = 12'b111111111111;
20'b00110000100100110100: color_data = 12'b111111111111;
20'b00110000100100110101: color_data = 12'b111111111111;
20'b00110000100100110110: color_data = 12'b111111111111;
20'b00110000100100110111: color_data = 12'b111111111111;
20'b00110000100100111000: color_data = 12'b111111111111;
20'b00110000100100111001: color_data = 12'b111111111111;
20'b00110000100100111010: color_data = 12'b111111111111;
20'b00110000100100111011: color_data = 12'b111111111111;
20'b00110000100100111100: color_data = 12'b111111111111;
20'b00110000100100111101: color_data = 12'b111111111111;
20'b00110000100100111110: color_data = 12'b111111111111;
20'b00110000100100111111: color_data = 12'b111111111111;
20'b00110000100101000100: color_data = 12'b111111111111;
20'b00110000100101000101: color_data = 12'b111111111111;
20'b00110000100101000110: color_data = 12'b111111111111;
20'b00110000100101000111: color_data = 12'b111111111111;
20'b00110000100101010000: color_data = 12'b111111111111;
20'b00110000100101010001: color_data = 12'b111111111111;
20'b00110000100101010010: color_data = 12'b111111111111;
20'b00110000100101010011: color_data = 12'b111111111111;
20'b00110000100101011000: color_data = 12'b111111111111;
20'b00110000100101011001: color_data = 12'b111111111111;
20'b00110000100101011010: color_data = 12'b111111111111;
20'b00110000100101011011: color_data = 12'b111111111111;
20'b00110000100101011100: color_data = 12'b111111111111;
20'b00110000100101011101: color_data = 12'b111111111111;
20'b00110000100101011110: color_data = 12'b111111111111;
20'b00110000100101011111: color_data = 12'b111111111111;
20'b00110000100101100000: color_data = 12'b111111111111;
20'b00110000100101100001: color_data = 12'b111111111111;
20'b00110000100101100010: color_data = 12'b111111111111;
20'b00110000100101100011: color_data = 12'b111111111111;
20'b00110000100101100100: color_data = 12'b111111111111;
20'b00110000100101100101: color_data = 12'b111111111111;
20'b00110000100101100110: color_data = 12'b111111111111;
20'b00110000100101100111: color_data = 12'b111111111111;
20'b00110000100101101100: color_data = 12'b111111111111;
20'b00110000100101101101: color_data = 12'b111111111111;
20'b00110000100101101110: color_data = 12'b111111111111;
20'b00110000100101101111: color_data = 12'b111111111111;
20'b00110000100110000100: color_data = 12'b111111111111;
20'b00110000100110000101: color_data = 12'b111111111111;
20'b00110000100110000110: color_data = 12'b111111111111;
20'b00110000100110000111: color_data = 12'b111111111111;
20'b00110000110100011100: color_data = 12'b111111111111;
20'b00110000110100011101: color_data = 12'b111111111111;
20'b00110000110100011110: color_data = 12'b111111111111;
20'b00110000110100011111: color_data = 12'b111111111111;
20'b00110000110100110000: color_data = 12'b111111111111;
20'b00110000110100110001: color_data = 12'b111111111111;
20'b00110000110100110010: color_data = 12'b111111111111;
20'b00110000110100110011: color_data = 12'b111111111111;
20'b00110000110100110100: color_data = 12'b111111111111;
20'b00110000110100110101: color_data = 12'b111111111111;
20'b00110000110100110110: color_data = 12'b111111111111;
20'b00110000110100110111: color_data = 12'b111111111111;
20'b00110000110100111000: color_data = 12'b111111111111;
20'b00110000110100111001: color_data = 12'b111111111111;
20'b00110000110100111010: color_data = 12'b111111111111;
20'b00110000110100111011: color_data = 12'b111111111111;
20'b00110000110100111100: color_data = 12'b111111111111;
20'b00110000110100111101: color_data = 12'b111111111111;
20'b00110000110100111110: color_data = 12'b111111111111;
20'b00110000110100111111: color_data = 12'b111111111111;
20'b00110000110101000100: color_data = 12'b111111111111;
20'b00110000110101000101: color_data = 12'b111111111111;
20'b00110000110101000110: color_data = 12'b111111111111;
20'b00110000110101000111: color_data = 12'b111111111111;
20'b00110000110101010000: color_data = 12'b111111111111;
20'b00110000110101010001: color_data = 12'b111111111111;
20'b00110000110101010010: color_data = 12'b111111111111;
20'b00110000110101010011: color_data = 12'b111111111111;
20'b00110000110101011000: color_data = 12'b111111111111;
20'b00110000110101011001: color_data = 12'b111111111111;
20'b00110000110101011010: color_data = 12'b111111111111;
20'b00110000110101011011: color_data = 12'b111111111111;
20'b00110000110101011100: color_data = 12'b111111111111;
20'b00110000110101011101: color_data = 12'b111111111111;
20'b00110000110101011110: color_data = 12'b111111111111;
20'b00110000110101011111: color_data = 12'b111111111111;
20'b00110000110101100000: color_data = 12'b111111111111;
20'b00110000110101100001: color_data = 12'b111111111111;
20'b00110000110101100010: color_data = 12'b111111111111;
20'b00110000110101100011: color_data = 12'b111111111111;
20'b00110000110101100100: color_data = 12'b111111111111;
20'b00110000110101100101: color_data = 12'b111111111111;
20'b00110000110101100110: color_data = 12'b111111111111;
20'b00110000110101100111: color_data = 12'b111111111111;
20'b00110000110101101100: color_data = 12'b111111111111;
20'b00110000110101101101: color_data = 12'b111111111111;
20'b00110000110101101110: color_data = 12'b111111111111;
20'b00110000110101101111: color_data = 12'b111111111111;
20'b00110000110110000100: color_data = 12'b111111111111;
20'b00110000110110000101: color_data = 12'b111111111111;
20'b00110000110110000110: color_data = 12'b111111111111;
20'b00110000110110000111: color_data = 12'b111111111111;
20'b00110001000100011100: color_data = 12'b111111111111;
20'b00110001000100011101: color_data = 12'b111111111111;
20'b00110001000100011110: color_data = 12'b111111111111;
20'b00110001000100011111: color_data = 12'b111111111111;
20'b00110001000100110000: color_data = 12'b111111111111;
20'b00110001000100110001: color_data = 12'b111111111111;
20'b00110001000100110010: color_data = 12'b111111111111;
20'b00110001000100110011: color_data = 12'b111111111111;
20'b00110001000100110100: color_data = 12'b111111111111;
20'b00110001000100110101: color_data = 12'b111111111111;
20'b00110001000100110110: color_data = 12'b111111111111;
20'b00110001000100110111: color_data = 12'b111111111111;
20'b00110001000100111000: color_data = 12'b111111111111;
20'b00110001000100111001: color_data = 12'b111111111111;
20'b00110001000100111010: color_data = 12'b111111111111;
20'b00110001000100111011: color_data = 12'b111111111111;
20'b00110001000100111100: color_data = 12'b111111111111;
20'b00110001000100111101: color_data = 12'b111111111111;
20'b00110001000100111110: color_data = 12'b111111111111;
20'b00110001000100111111: color_data = 12'b111111111111;
20'b00110001000101000100: color_data = 12'b111111111111;
20'b00110001000101000101: color_data = 12'b111111111111;
20'b00110001000101000110: color_data = 12'b111111111111;
20'b00110001000101000111: color_data = 12'b111111111111;
20'b00110001000101010000: color_data = 12'b111111111111;
20'b00110001000101010001: color_data = 12'b111111111111;
20'b00110001000101010010: color_data = 12'b111111111111;
20'b00110001000101010011: color_data = 12'b111111111111;
20'b00110001000101011000: color_data = 12'b111111111111;
20'b00110001000101011001: color_data = 12'b111111111111;
20'b00110001000101011010: color_data = 12'b111111111111;
20'b00110001000101011011: color_data = 12'b111111111111;
20'b00110001000101011100: color_data = 12'b111111111111;
20'b00110001000101011101: color_data = 12'b111111111111;
20'b00110001000101011110: color_data = 12'b111111111111;
20'b00110001000101011111: color_data = 12'b111111111111;
20'b00110001000101100000: color_data = 12'b111111111111;
20'b00110001000101100001: color_data = 12'b111111111111;
20'b00110001000101100010: color_data = 12'b111111111111;
20'b00110001000101100011: color_data = 12'b111111111111;
20'b00110001000101100100: color_data = 12'b111111111111;
20'b00110001000101100101: color_data = 12'b111111111111;
20'b00110001000101100110: color_data = 12'b111111111111;
20'b00110001000101100111: color_data = 12'b111111111111;
20'b00110001000101101100: color_data = 12'b111111111111;
20'b00110001000101101101: color_data = 12'b111111111111;
20'b00110001000101101110: color_data = 12'b111111111111;
20'b00110001000101101111: color_data = 12'b111111111111;
20'b00110001000110000100: color_data = 12'b111111111111;
20'b00110001000110000101: color_data = 12'b111111111111;
20'b00110001000110000110: color_data = 12'b111111111111;
20'b00110001000110000111: color_data = 12'b111111111111;
20'b00110001010100011100: color_data = 12'b111111111111;
20'b00110001010100011101: color_data = 12'b111111111111;
20'b00110001010100011110: color_data = 12'b111111111111;
20'b00110001010100011111: color_data = 12'b111111111111;
20'b00110001010100110000: color_data = 12'b111111111111;
20'b00110001010100110001: color_data = 12'b111111111111;
20'b00110001010100110010: color_data = 12'b111111111111;
20'b00110001010100110011: color_data = 12'b111111111111;
20'b00110001010101000100: color_data = 12'b111111111111;
20'b00110001010101000101: color_data = 12'b111111111111;
20'b00110001010101000110: color_data = 12'b111111111111;
20'b00110001010101000111: color_data = 12'b111111111111;
20'b00110001010101010000: color_data = 12'b111111111111;
20'b00110001010101010001: color_data = 12'b111111111111;
20'b00110001010101010010: color_data = 12'b111111111111;
20'b00110001010101010011: color_data = 12'b111111111111;
20'b00110001010101011000: color_data = 12'b111111111111;
20'b00110001010101011001: color_data = 12'b111111111111;
20'b00110001010101011010: color_data = 12'b111111111111;
20'b00110001010101011011: color_data = 12'b111111111111;
20'b00110001010101101100: color_data = 12'b111111111111;
20'b00110001010101101101: color_data = 12'b111111111111;
20'b00110001010101101110: color_data = 12'b111111111111;
20'b00110001010101101111: color_data = 12'b111111111111;
20'b00110001010110000100: color_data = 12'b111111111111;
20'b00110001010110000101: color_data = 12'b111111111111;
20'b00110001010110000110: color_data = 12'b111111111111;
20'b00110001010110000111: color_data = 12'b111111111111;
20'b00110001100100011100: color_data = 12'b111111111111;
20'b00110001100100011101: color_data = 12'b111111111111;
20'b00110001100100011110: color_data = 12'b111111111111;
20'b00110001100100011111: color_data = 12'b111111111111;
20'b00110001100100110000: color_data = 12'b111111111111;
20'b00110001100100110001: color_data = 12'b111111111111;
20'b00110001100100110010: color_data = 12'b111111111111;
20'b00110001100100110011: color_data = 12'b111111111111;
20'b00110001100101000100: color_data = 12'b111111111111;
20'b00110001100101000101: color_data = 12'b111111111111;
20'b00110001100101000110: color_data = 12'b111111111111;
20'b00110001100101000111: color_data = 12'b111111111111;
20'b00110001100101010000: color_data = 12'b111111111111;
20'b00110001100101010001: color_data = 12'b111111111111;
20'b00110001100101010010: color_data = 12'b111111111111;
20'b00110001100101010011: color_data = 12'b111111111111;
20'b00110001100101011000: color_data = 12'b111111111111;
20'b00110001100101011001: color_data = 12'b111111111111;
20'b00110001100101011010: color_data = 12'b111111111111;
20'b00110001100101011011: color_data = 12'b111111111111;
20'b00110001100101101100: color_data = 12'b111111111111;
20'b00110001100101101101: color_data = 12'b111111111111;
20'b00110001100101101110: color_data = 12'b111111111111;
20'b00110001100101101111: color_data = 12'b111111111111;
20'b00110001100110000100: color_data = 12'b111111111111;
20'b00110001100110000101: color_data = 12'b111111111111;
20'b00110001100110000110: color_data = 12'b111111111111;
20'b00110001100110000111: color_data = 12'b111111111111;
20'b00110001110100011100: color_data = 12'b111111111111;
20'b00110001110100011101: color_data = 12'b111111111111;
20'b00110001110100011110: color_data = 12'b111111111111;
20'b00110001110100011111: color_data = 12'b111111111111;
20'b00110001110100110000: color_data = 12'b111111111111;
20'b00110001110100110001: color_data = 12'b111111111111;
20'b00110001110100110010: color_data = 12'b111111111111;
20'b00110001110100110011: color_data = 12'b111111111111;
20'b00110001110101000100: color_data = 12'b111111111111;
20'b00110001110101000101: color_data = 12'b111111111111;
20'b00110001110101000110: color_data = 12'b111111111111;
20'b00110001110101000111: color_data = 12'b111111111111;
20'b00110001110101010000: color_data = 12'b111111111111;
20'b00110001110101010001: color_data = 12'b111111111111;
20'b00110001110101010010: color_data = 12'b111111111111;
20'b00110001110101010011: color_data = 12'b111111111111;
20'b00110001110101011000: color_data = 12'b111111111111;
20'b00110001110101011001: color_data = 12'b111111111111;
20'b00110001110101011010: color_data = 12'b111111111111;
20'b00110001110101011011: color_data = 12'b111111111111;
20'b00110001110101101100: color_data = 12'b111111111111;
20'b00110001110101101101: color_data = 12'b111111111111;
20'b00110001110101101110: color_data = 12'b111111111111;
20'b00110001110101101111: color_data = 12'b111111111111;
20'b00110001110110000100: color_data = 12'b111111111111;
20'b00110001110110000101: color_data = 12'b111111111111;
20'b00110001110110000110: color_data = 12'b111111111111;
20'b00110001110110000111: color_data = 12'b111111111111;
20'b00110010000100010101: color_data = 12'b111111111111;
20'b00110010000100010110: color_data = 12'b111111111111;
20'b00110010000100010111: color_data = 12'b111111111111;
20'b00110010000100011000: color_data = 12'b111111111111;
20'b00110010000100011100: color_data = 12'b111111111111;
20'b00110010000100011101: color_data = 12'b111111111111;
20'b00110010000100011110: color_data = 12'b111111111111;
20'b00110010000100011111: color_data = 12'b111111111111;
20'b00110010000100110000: color_data = 12'b111111111111;
20'b00110010000100110001: color_data = 12'b111111111111;
20'b00110010000100110010: color_data = 12'b111111111111;
20'b00110010000100110011: color_data = 12'b111111111111;
20'b00110010000100110100: color_data = 12'b111111111111;
20'b00110010000100110101: color_data = 12'b111111111111;
20'b00110010000100110110: color_data = 12'b111111111111;
20'b00110010000100110111: color_data = 12'b111111111111;
20'b00110010000100111000: color_data = 12'b111111111111;
20'b00110010000100111001: color_data = 12'b111111111111;
20'b00110010000100111010: color_data = 12'b111111111111;
20'b00110010000100111011: color_data = 12'b111111111111;
20'b00110010000100111100: color_data = 12'b111111111111;
20'b00110010000100111101: color_data = 12'b111111111111;
20'b00110010000100111110: color_data = 12'b111111111111;
20'b00110010000100111111: color_data = 12'b111111111111;
20'b00110010000101000100: color_data = 12'b111111111111;
20'b00110010000101000101: color_data = 12'b111111111111;
20'b00110010000101000110: color_data = 12'b111111111111;
20'b00110010000101000111: color_data = 12'b111111111111;
20'b00110010000101010000: color_data = 12'b111111111111;
20'b00110010000101010001: color_data = 12'b111111111111;
20'b00110010000101010010: color_data = 12'b111111111111;
20'b00110010000101010011: color_data = 12'b111111111111;
20'b00110010000101011000: color_data = 12'b111111111111;
20'b00110010000101011001: color_data = 12'b111111111111;
20'b00110010000101011010: color_data = 12'b111111111111;
20'b00110010000101011011: color_data = 12'b111111111111;
20'b00110010000101011100: color_data = 12'b111111111111;
20'b00110010000101011101: color_data = 12'b111111111111;
20'b00110010000101011110: color_data = 12'b111111111111;
20'b00110010000101011111: color_data = 12'b111111111111;
20'b00110010000101100000: color_data = 12'b111111111111;
20'b00110010000101100001: color_data = 12'b111111111111;
20'b00110010000101100010: color_data = 12'b111111111111;
20'b00110010000101100011: color_data = 12'b111111111111;
20'b00110010000101100100: color_data = 12'b111111111111;
20'b00110010000101100101: color_data = 12'b111111111111;
20'b00110010000101100110: color_data = 12'b111111111111;
20'b00110010000101100111: color_data = 12'b111111111111;
20'b00110010000101101100: color_data = 12'b111111111111;
20'b00110010000101101101: color_data = 12'b111111111111;
20'b00110010000101101110: color_data = 12'b111111111111;
20'b00110010000101101111: color_data = 12'b111111111111;
20'b00110010000110000100: color_data = 12'b111111111111;
20'b00110010000110000101: color_data = 12'b111111111111;
20'b00110010000110000110: color_data = 12'b111111111111;
20'b00110010000110000111: color_data = 12'b111111111111;
20'b00110010010100010101: color_data = 12'b111111111111;
20'b00110010010100010110: color_data = 12'b111111111111;
20'b00110010010100010111: color_data = 12'b111111111111;
20'b00110010010100011000: color_data = 12'b111111111111;
20'b00110010010100011100: color_data = 12'b111111111111;
20'b00110010010100011101: color_data = 12'b111111111111;
20'b00110010010100011110: color_data = 12'b111111111111;
20'b00110010010100011111: color_data = 12'b111111111111;
20'b00110010010100110000: color_data = 12'b111111111111;
20'b00110010010100110001: color_data = 12'b111111111111;
20'b00110010010100110010: color_data = 12'b111111111111;
20'b00110010010100110011: color_data = 12'b111111111111;
20'b00110010010100110100: color_data = 12'b111111111111;
20'b00110010010100110101: color_data = 12'b111111111111;
20'b00110010010100110110: color_data = 12'b111111111111;
20'b00110010010100110111: color_data = 12'b111111111111;
20'b00110010010100111000: color_data = 12'b111111111111;
20'b00110010010100111001: color_data = 12'b111111111111;
20'b00110010010100111010: color_data = 12'b111111111111;
20'b00110010010100111011: color_data = 12'b111111111111;
20'b00110010010100111100: color_data = 12'b111111111111;
20'b00110010010100111101: color_data = 12'b111111111111;
20'b00110010010100111110: color_data = 12'b111111111111;
20'b00110010010100111111: color_data = 12'b111111111111;
20'b00110010010101000100: color_data = 12'b111111111111;
20'b00110010010101000101: color_data = 12'b111111111111;
20'b00110010010101000110: color_data = 12'b111111111111;
20'b00110010010101000111: color_data = 12'b111111111111;
20'b00110010010101010000: color_data = 12'b111111111111;
20'b00110010010101010001: color_data = 12'b111111111111;
20'b00110010010101010010: color_data = 12'b111111111111;
20'b00110010010101010011: color_data = 12'b111111111111;
20'b00110010010101011000: color_data = 12'b111111111111;
20'b00110010010101011001: color_data = 12'b111111111111;
20'b00110010010101011010: color_data = 12'b111111111111;
20'b00110010010101011011: color_data = 12'b111111111111;
20'b00110010010101011100: color_data = 12'b111111111111;
20'b00110010010101011101: color_data = 12'b111111111111;
20'b00110010010101011110: color_data = 12'b111111111111;
20'b00110010010101011111: color_data = 12'b111111111111;
20'b00110010010101100000: color_data = 12'b111111111111;
20'b00110010010101100001: color_data = 12'b111111111111;
20'b00110010010101100010: color_data = 12'b111111111111;
20'b00110010010101100011: color_data = 12'b111111111111;
20'b00110010010101100100: color_data = 12'b111111111111;
20'b00110010010101100101: color_data = 12'b111111111111;
20'b00110010010101100110: color_data = 12'b111111111111;
20'b00110010010101100111: color_data = 12'b111111111111;
20'b00110010010101101100: color_data = 12'b111111111111;
20'b00110010010101101101: color_data = 12'b111111111111;
20'b00110010010101101110: color_data = 12'b111111111111;
20'b00110010010101101111: color_data = 12'b111111111111;
20'b00110010010110000100: color_data = 12'b111111111111;
20'b00110010010110000101: color_data = 12'b111111111111;
20'b00110010010110000110: color_data = 12'b111111111111;
20'b00110010010110000111: color_data = 12'b111111111111;
20'b00110010100100010101: color_data = 12'b111111111111;
20'b00110010100100010110: color_data = 12'b111111111111;
20'b00110010100100010111: color_data = 12'b111111111111;
20'b00110010100100011000: color_data = 12'b111111111111;
20'b00110010100100011100: color_data = 12'b111111111111;
20'b00110010100100011101: color_data = 12'b111111111111;
20'b00110010100100011110: color_data = 12'b111111111111;
20'b00110010100100011111: color_data = 12'b111111111111;
20'b00110010100100110000: color_data = 12'b111111111111;
20'b00110010100100110001: color_data = 12'b111111111111;
20'b00110010100100110010: color_data = 12'b111111111111;
20'b00110010100100110011: color_data = 12'b111111111111;
20'b00110010100100110100: color_data = 12'b111111111111;
20'b00110010100100110101: color_data = 12'b111111111111;
20'b00110010100100110110: color_data = 12'b111111111111;
20'b00110010100100110111: color_data = 12'b111111111111;
20'b00110010100100111000: color_data = 12'b111111111111;
20'b00110010100100111001: color_data = 12'b111111111111;
20'b00110010100100111010: color_data = 12'b111111111111;
20'b00110010100100111011: color_data = 12'b111111111111;
20'b00110010100100111100: color_data = 12'b111111111111;
20'b00110010100100111101: color_data = 12'b111111111111;
20'b00110010100100111110: color_data = 12'b111111111111;
20'b00110010100100111111: color_data = 12'b111111111111;
20'b00110010100101000100: color_data = 12'b111111111111;
20'b00110010100101000101: color_data = 12'b111111111111;
20'b00110010100101000110: color_data = 12'b111111111111;
20'b00110010100101000111: color_data = 12'b111111111111;
20'b00110010100101010000: color_data = 12'b111111111111;
20'b00110010100101010001: color_data = 12'b111111111111;
20'b00110010100101010010: color_data = 12'b111111111111;
20'b00110010100101010011: color_data = 12'b111111111111;
20'b00110010100101011000: color_data = 12'b111111111111;
20'b00110010100101011001: color_data = 12'b111111111111;
20'b00110010100101011010: color_data = 12'b111111111111;
20'b00110010100101011011: color_data = 12'b111111111111;
20'b00110010100101011100: color_data = 12'b111111111111;
20'b00110010100101011101: color_data = 12'b111111111111;
20'b00110010100101011110: color_data = 12'b111111111111;
20'b00110010100101011111: color_data = 12'b111111111111;
20'b00110010100101100000: color_data = 12'b111111111111;
20'b00110010100101100001: color_data = 12'b111111111111;
20'b00110010100101100010: color_data = 12'b111111111111;
20'b00110010100101100011: color_data = 12'b111111111111;
20'b00110010100101100100: color_data = 12'b111111111111;
20'b00110010100101100101: color_data = 12'b111111111111;
20'b00110010100101100110: color_data = 12'b111111111111;
20'b00110010100101100111: color_data = 12'b111111111111;
20'b00110010100101101100: color_data = 12'b111111111111;
20'b00110010100101101101: color_data = 12'b111111111111;
20'b00110010100101101110: color_data = 12'b111111111111;
20'b00110010100101101111: color_data = 12'b111111111111;
20'b00110010100110000100: color_data = 12'b111111111111;
20'b00110010100110000101: color_data = 12'b111111111111;
20'b00110010100110000110: color_data = 12'b111111111111;
20'b00110010100110000111: color_data = 12'b111111111111;
20'b00110010110100010101: color_data = 12'b111111111111;
20'b00110010110100010110: color_data = 12'b111111111111;
20'b00110010110100010111: color_data = 12'b111111111111;
20'b00110010110100011000: color_data = 12'b111111111111;
20'b00110010110100011100: color_data = 12'b111111111111;
20'b00110010110100011101: color_data = 12'b111111111111;
20'b00110010110100011110: color_data = 12'b111111111111;
20'b00110010110100011111: color_data = 12'b111111111111;
20'b00110010110100110000: color_data = 12'b111111111111;
20'b00110010110100110001: color_data = 12'b111111111111;
20'b00110010110100110010: color_data = 12'b111111111111;
20'b00110010110100110011: color_data = 12'b111111111111;
20'b00110010110100110100: color_data = 12'b111111111111;
20'b00110010110100110101: color_data = 12'b111111111111;
20'b00110010110100110110: color_data = 12'b111111111111;
20'b00110010110100110111: color_data = 12'b111111111111;
20'b00110010110100111000: color_data = 12'b111111111111;
20'b00110010110100111001: color_data = 12'b111111111111;
20'b00110010110100111010: color_data = 12'b111111111111;
20'b00110010110100111011: color_data = 12'b111111111111;
20'b00110010110100111100: color_data = 12'b111111111111;
20'b00110010110100111101: color_data = 12'b111111111111;
20'b00110010110100111110: color_data = 12'b111111111111;
20'b00110010110100111111: color_data = 12'b111111111111;
20'b00110010110101000100: color_data = 12'b111111111111;
20'b00110010110101000101: color_data = 12'b111111111111;
20'b00110010110101000110: color_data = 12'b111111111111;
20'b00110010110101000111: color_data = 12'b111111111111;
20'b00110010110101010000: color_data = 12'b111111111111;
20'b00110010110101010001: color_data = 12'b111111111111;
20'b00110010110101010010: color_data = 12'b111111111111;
20'b00110010110101010011: color_data = 12'b111111111111;
20'b00110010110101011000: color_data = 12'b111111111111;
20'b00110010110101011001: color_data = 12'b111111111111;
20'b00110010110101011010: color_data = 12'b111111111111;
20'b00110010110101011011: color_data = 12'b111111111111;
20'b00110010110101011100: color_data = 12'b111111111111;
20'b00110010110101011101: color_data = 12'b111111111111;
20'b00110010110101011110: color_data = 12'b111111111111;
20'b00110010110101011111: color_data = 12'b111111111111;
20'b00110010110101100000: color_data = 12'b111111111111;
20'b00110010110101100001: color_data = 12'b111111111111;
20'b00110010110101100010: color_data = 12'b111111111111;
20'b00110010110101100011: color_data = 12'b111111111111;
20'b00110010110101100100: color_data = 12'b111111111111;
20'b00110010110101100101: color_data = 12'b111111111111;
20'b00110010110101100110: color_data = 12'b111111111111;
20'b00110010110101100111: color_data = 12'b111111111111;
20'b00110010110101101100: color_data = 12'b111111111111;
20'b00110010110101101101: color_data = 12'b111111111111;
20'b00110010110101101110: color_data = 12'b111111111111;
20'b00110010110101101111: color_data = 12'b111111111111;
20'b00110010110110000100: color_data = 12'b111111111111;
20'b00110010110110000101: color_data = 12'b111111111111;
20'b00110010110110000110: color_data = 12'b111111111111;
20'b00110010110110000111: color_data = 12'b111111111111;
20'b00110011000100011100: color_data = 12'b111111111111;
20'b00110011000100011101: color_data = 12'b111111111111;
20'b00110011000100011110: color_data = 12'b111111111111;
20'b00110011000100011111: color_data = 12'b111111111111;
20'b00110011000100110000: color_data = 12'b111111111111;
20'b00110011000100110001: color_data = 12'b111111111111;
20'b00110011000100110010: color_data = 12'b111111111111;
20'b00110011000100110011: color_data = 12'b111111111111;
20'b00110011000101000100: color_data = 12'b111111111111;
20'b00110011000101000101: color_data = 12'b111111111111;
20'b00110011000101000110: color_data = 12'b111111111111;
20'b00110011000101000111: color_data = 12'b111111111111;
20'b00110011000101010000: color_data = 12'b111111111111;
20'b00110011000101010001: color_data = 12'b111111111111;
20'b00110011000101010010: color_data = 12'b111111111111;
20'b00110011000101010011: color_data = 12'b111111111111;
20'b00110011000101011000: color_data = 12'b111111111111;
20'b00110011000101011001: color_data = 12'b111111111111;
20'b00110011000101011010: color_data = 12'b111111111111;
20'b00110011000101011011: color_data = 12'b111111111111;
20'b00110011000101101100: color_data = 12'b111111111111;
20'b00110011000101101101: color_data = 12'b111111111111;
20'b00110011000101101110: color_data = 12'b111111111111;
20'b00110011000101101111: color_data = 12'b111111111111;
20'b00110011000110000100: color_data = 12'b111111111111;
20'b00110011000110000101: color_data = 12'b111111111111;
20'b00110011000110000110: color_data = 12'b111111111111;
20'b00110011000110000111: color_data = 12'b111111111111;
20'b00110011010100011100: color_data = 12'b111111111111;
20'b00110011010100011101: color_data = 12'b111111111111;
20'b00110011010100011110: color_data = 12'b111111111111;
20'b00110011010100011111: color_data = 12'b111111111111;
20'b00110011010100110000: color_data = 12'b111111111111;
20'b00110011010100110001: color_data = 12'b111111111111;
20'b00110011010100110010: color_data = 12'b111111111111;
20'b00110011010100110011: color_data = 12'b111111111111;
20'b00110011010101000100: color_data = 12'b111111111111;
20'b00110011010101000101: color_data = 12'b111111111111;
20'b00110011010101000110: color_data = 12'b111111111111;
20'b00110011010101000111: color_data = 12'b111111111111;
20'b00110011010101010000: color_data = 12'b111111111111;
20'b00110011010101010001: color_data = 12'b111111111111;
20'b00110011010101010010: color_data = 12'b111111111111;
20'b00110011010101010011: color_data = 12'b111111111111;
20'b00110011010101011000: color_data = 12'b111111111111;
20'b00110011010101011001: color_data = 12'b111111111111;
20'b00110011010101011010: color_data = 12'b111111111111;
20'b00110011010101011011: color_data = 12'b111111111111;
20'b00110011010101101100: color_data = 12'b111111111111;
20'b00110011010101101101: color_data = 12'b111111111111;
20'b00110011010101101110: color_data = 12'b111111111111;
20'b00110011010101101111: color_data = 12'b111111111111;
20'b00110011010110000100: color_data = 12'b111111111111;
20'b00110011010110000101: color_data = 12'b111111111111;
20'b00110011010110000110: color_data = 12'b111111111111;
20'b00110011010110000111: color_data = 12'b111111111111;
20'b00110011100100011100: color_data = 12'b111111111111;
20'b00110011100100011101: color_data = 12'b111111111111;
20'b00110011100100011110: color_data = 12'b111111111111;
20'b00110011100100011111: color_data = 12'b111111111111;
20'b00110011100100110000: color_data = 12'b111111111111;
20'b00110011100100110001: color_data = 12'b111111111111;
20'b00110011100100110010: color_data = 12'b111111111111;
20'b00110011100100110011: color_data = 12'b111111111111;
20'b00110011100101000100: color_data = 12'b111111111111;
20'b00110011100101000101: color_data = 12'b111111111111;
20'b00110011100101000110: color_data = 12'b111111111111;
20'b00110011100101000111: color_data = 12'b111111111111;
20'b00110011100101010000: color_data = 12'b111111111111;
20'b00110011100101010001: color_data = 12'b111111111111;
20'b00110011100101010010: color_data = 12'b111111111111;
20'b00110011100101010011: color_data = 12'b111111111111;
20'b00110011100101011000: color_data = 12'b111111111111;
20'b00110011100101011001: color_data = 12'b111111111111;
20'b00110011100101011010: color_data = 12'b111111111111;
20'b00110011100101011011: color_data = 12'b111111111111;
20'b00110011100101101100: color_data = 12'b111111111111;
20'b00110011100101101101: color_data = 12'b111111111111;
20'b00110011100101101110: color_data = 12'b111111111111;
20'b00110011100101101111: color_data = 12'b111111111111;
20'b00110011100110000100: color_data = 12'b111111111111;
20'b00110011100110000101: color_data = 12'b111111111111;
20'b00110011100110000110: color_data = 12'b111111111111;
20'b00110011100110000111: color_data = 12'b111111111111;
20'b00110011110100011100: color_data = 12'b111111111111;
20'b00110011110100011101: color_data = 12'b111111111111;
20'b00110011110100011110: color_data = 12'b111111111111;
20'b00110011110100011111: color_data = 12'b111111111111;
20'b00110011110100100000: color_data = 12'b111111111111;
20'b00110011110100100001: color_data = 12'b111111111111;
20'b00110011110100100010: color_data = 12'b111111111111;
20'b00110011110100100011: color_data = 12'b111111111111;
20'b00110011110100100100: color_data = 12'b111111111111;
20'b00110011110100100101: color_data = 12'b111111111111;
20'b00110011110100100110: color_data = 12'b111111111111;
20'b00110011110100100111: color_data = 12'b111111111111;
20'b00110011110100101000: color_data = 12'b111111111111;
20'b00110011110100101001: color_data = 12'b111111111111;
20'b00110011110100101010: color_data = 12'b111111111111;
20'b00110011110100101011: color_data = 12'b111111111111;
20'b00110011110100110000: color_data = 12'b111111111111;
20'b00110011110100110001: color_data = 12'b111111111111;
20'b00110011110100110010: color_data = 12'b111111111111;
20'b00110011110100110011: color_data = 12'b111111111111;
20'b00110011110100110100: color_data = 12'b111111111111;
20'b00110011110100110101: color_data = 12'b111111111111;
20'b00110011110100110110: color_data = 12'b111111111111;
20'b00110011110100110111: color_data = 12'b111111111111;
20'b00110011110100111000: color_data = 12'b111111111111;
20'b00110011110100111001: color_data = 12'b111111111111;
20'b00110011110100111010: color_data = 12'b111111111111;
20'b00110011110100111011: color_data = 12'b111111111111;
20'b00110011110100111100: color_data = 12'b111111111111;
20'b00110011110100111101: color_data = 12'b111111111111;
20'b00110011110100111110: color_data = 12'b111111111111;
20'b00110011110100111111: color_data = 12'b111111111111;
20'b00110011110101000100: color_data = 12'b111111111111;
20'b00110011110101000101: color_data = 12'b111111111111;
20'b00110011110101000110: color_data = 12'b111111111111;
20'b00110011110101000111: color_data = 12'b111111111111;
20'b00110011110101001000: color_data = 12'b111111111111;
20'b00110011110101001001: color_data = 12'b111111111111;
20'b00110011110101001010: color_data = 12'b111111111111;
20'b00110011110101001011: color_data = 12'b111111111111;
20'b00110011110101001100: color_data = 12'b111111111111;
20'b00110011110101001101: color_data = 12'b111111111111;
20'b00110011110101001110: color_data = 12'b111111111111;
20'b00110011110101001111: color_data = 12'b111111111111;
20'b00110011110101011000: color_data = 12'b111111111111;
20'b00110011110101011001: color_data = 12'b111111111111;
20'b00110011110101011010: color_data = 12'b111111111111;
20'b00110011110101011011: color_data = 12'b111111111111;
20'b00110011110101011100: color_data = 12'b111111111111;
20'b00110011110101011101: color_data = 12'b111111111111;
20'b00110011110101011110: color_data = 12'b111111111111;
20'b00110011110101011111: color_data = 12'b111111111111;
20'b00110011110101100000: color_data = 12'b111111111111;
20'b00110011110101100001: color_data = 12'b111111111111;
20'b00110011110101100010: color_data = 12'b111111111111;
20'b00110011110101100011: color_data = 12'b111111111111;
20'b00110011110101100100: color_data = 12'b111111111111;
20'b00110011110101100101: color_data = 12'b111111111111;
20'b00110011110101100110: color_data = 12'b111111111111;
20'b00110011110101100111: color_data = 12'b111111111111;
20'b00110011110101101100: color_data = 12'b111111111111;
20'b00110011110101101101: color_data = 12'b111111111111;
20'b00110011110101101110: color_data = 12'b111111111111;
20'b00110011110101101111: color_data = 12'b111111111111;
20'b00110011110101110000: color_data = 12'b111111111111;
20'b00110011110101110001: color_data = 12'b111111111111;
20'b00110011110101110010: color_data = 12'b111111111111;
20'b00110011110101110011: color_data = 12'b111111111111;
20'b00110011110101110100: color_data = 12'b111111111111;
20'b00110011110101110101: color_data = 12'b111111111111;
20'b00110011110101110110: color_data = 12'b111111111111;
20'b00110011110101110111: color_data = 12'b111111111111;
20'b00110011110101111000: color_data = 12'b111111111111;
20'b00110011110101111001: color_data = 12'b111111111111;
20'b00110011110101111010: color_data = 12'b111111111111;
20'b00110011110101111011: color_data = 12'b111111111111;
20'b00110011110110000100: color_data = 12'b111111111111;
20'b00110011110110000101: color_data = 12'b111111111111;
20'b00110011110110000110: color_data = 12'b111111111111;
20'b00110011110110000111: color_data = 12'b111111111111;
20'b00110100000100011100: color_data = 12'b111111111111;
20'b00110100000100011101: color_data = 12'b111111111111;
20'b00110100000100011110: color_data = 12'b111111111111;
20'b00110100000100011111: color_data = 12'b111111111111;
20'b00110100000100100000: color_data = 12'b111111111111;
20'b00110100000100100001: color_data = 12'b111111111111;
20'b00110100000100100010: color_data = 12'b111111111111;
20'b00110100000100100011: color_data = 12'b111111111111;
20'b00110100000100100100: color_data = 12'b111111111111;
20'b00110100000100100101: color_data = 12'b111111111111;
20'b00110100000100100110: color_data = 12'b111111111111;
20'b00110100000100100111: color_data = 12'b111111111111;
20'b00110100000100101000: color_data = 12'b111111111111;
20'b00110100000100101001: color_data = 12'b111111111111;
20'b00110100000100101010: color_data = 12'b111111111111;
20'b00110100000100101011: color_data = 12'b111111111111;
20'b00110100000100110000: color_data = 12'b111111111111;
20'b00110100000100110001: color_data = 12'b111111111111;
20'b00110100000100110010: color_data = 12'b111111111111;
20'b00110100000100110011: color_data = 12'b111111111111;
20'b00110100000100110100: color_data = 12'b111111111111;
20'b00110100000100110101: color_data = 12'b111111111111;
20'b00110100000100110110: color_data = 12'b111111111111;
20'b00110100000100110111: color_data = 12'b111111111111;
20'b00110100000100111000: color_data = 12'b111111111111;
20'b00110100000100111001: color_data = 12'b111111111111;
20'b00110100000100111010: color_data = 12'b111111111111;
20'b00110100000100111011: color_data = 12'b111111111111;
20'b00110100000100111100: color_data = 12'b111111111111;
20'b00110100000100111101: color_data = 12'b111111111111;
20'b00110100000100111110: color_data = 12'b111111111111;
20'b00110100000100111111: color_data = 12'b111111111111;
20'b00110100000101000100: color_data = 12'b111111111111;
20'b00110100000101000101: color_data = 12'b111111111111;
20'b00110100000101000110: color_data = 12'b111111111111;
20'b00110100000101000111: color_data = 12'b111111111111;
20'b00110100000101001000: color_data = 12'b111111111111;
20'b00110100000101001001: color_data = 12'b111111111111;
20'b00110100000101001010: color_data = 12'b111111111111;
20'b00110100000101001011: color_data = 12'b111111111111;
20'b00110100000101001100: color_data = 12'b111111111111;
20'b00110100000101001101: color_data = 12'b111111111111;
20'b00110100000101001110: color_data = 12'b111111111111;
20'b00110100000101001111: color_data = 12'b111111111111;
20'b00110100000101011000: color_data = 12'b111111111111;
20'b00110100000101011001: color_data = 12'b111111111111;
20'b00110100000101011010: color_data = 12'b111111111111;
20'b00110100000101011011: color_data = 12'b111111111111;
20'b00110100000101011100: color_data = 12'b111111111111;
20'b00110100000101011101: color_data = 12'b111111111111;
20'b00110100000101011110: color_data = 12'b111111111111;
20'b00110100000101011111: color_data = 12'b111111111111;
20'b00110100000101100000: color_data = 12'b111111111111;
20'b00110100000101100001: color_data = 12'b111111111111;
20'b00110100000101100010: color_data = 12'b111111111111;
20'b00110100000101100011: color_data = 12'b111111111111;
20'b00110100000101100100: color_data = 12'b111111111111;
20'b00110100000101100101: color_data = 12'b111111111111;
20'b00110100000101100110: color_data = 12'b111111111111;
20'b00110100000101100111: color_data = 12'b111111111111;
20'b00110100000101101100: color_data = 12'b111111111111;
20'b00110100000101101101: color_data = 12'b111111111111;
20'b00110100000101101110: color_data = 12'b111111111111;
20'b00110100000101101111: color_data = 12'b111111111111;
20'b00110100000101110000: color_data = 12'b111111111111;
20'b00110100000101110001: color_data = 12'b111111111111;
20'b00110100000101110010: color_data = 12'b111111111111;
20'b00110100000101110011: color_data = 12'b111111111111;
20'b00110100000101110100: color_data = 12'b111111111111;
20'b00110100000101110101: color_data = 12'b111111111111;
20'b00110100000101110110: color_data = 12'b111111111111;
20'b00110100000101110111: color_data = 12'b111111111111;
20'b00110100000101111000: color_data = 12'b111111111111;
20'b00110100000101111001: color_data = 12'b111111111111;
20'b00110100000101111010: color_data = 12'b111111111111;
20'b00110100000101111011: color_data = 12'b111111111111;
20'b00110100000110000100: color_data = 12'b111111111111;
20'b00110100000110000101: color_data = 12'b111111111111;
20'b00110100000110000110: color_data = 12'b111111111111;
20'b00110100000110000111: color_data = 12'b111111111111;
20'b00110100010100011100: color_data = 12'b111111111111;
20'b00110100010100011101: color_data = 12'b111111111111;
20'b00110100010100011110: color_data = 12'b111111111111;
20'b00110100010100011111: color_data = 12'b111111111111;
20'b00110100010100100000: color_data = 12'b111111111111;
20'b00110100010100100001: color_data = 12'b111111111111;
20'b00110100010100100010: color_data = 12'b111111111111;
20'b00110100010100100011: color_data = 12'b111111111111;
20'b00110100010100100100: color_data = 12'b111111111111;
20'b00110100010100100101: color_data = 12'b111111111111;
20'b00110100010100100110: color_data = 12'b111111111111;
20'b00110100010100100111: color_data = 12'b111111111111;
20'b00110100010100101000: color_data = 12'b111111111111;
20'b00110100010100101001: color_data = 12'b111111111111;
20'b00110100010100101010: color_data = 12'b111111111111;
20'b00110100010100101011: color_data = 12'b111111111111;
20'b00110100010100110000: color_data = 12'b111111111111;
20'b00110100010100110001: color_data = 12'b111111111111;
20'b00110100010100110010: color_data = 12'b111111111111;
20'b00110100010100110011: color_data = 12'b111111111111;
20'b00110100010100110100: color_data = 12'b111111111111;
20'b00110100010100110101: color_data = 12'b111111111111;
20'b00110100010100110110: color_data = 12'b111111111111;
20'b00110100010100110111: color_data = 12'b111111111111;
20'b00110100010100111000: color_data = 12'b111111111111;
20'b00110100010100111001: color_data = 12'b111111111111;
20'b00110100010100111010: color_data = 12'b111111111111;
20'b00110100010100111011: color_data = 12'b111111111111;
20'b00110100010100111100: color_data = 12'b111111111111;
20'b00110100010100111101: color_data = 12'b111111111111;
20'b00110100010100111110: color_data = 12'b111111111111;
20'b00110100010100111111: color_data = 12'b111111111111;
20'b00110100010101000100: color_data = 12'b111111111111;
20'b00110100010101000101: color_data = 12'b111111111111;
20'b00110100010101000110: color_data = 12'b111111111111;
20'b00110100010101000111: color_data = 12'b111111111111;
20'b00110100010101001000: color_data = 12'b111111111111;
20'b00110100010101001001: color_data = 12'b111111111111;
20'b00110100010101001010: color_data = 12'b111111111111;
20'b00110100010101001011: color_data = 12'b111111111111;
20'b00110100010101001100: color_data = 12'b111111111111;
20'b00110100010101001101: color_data = 12'b111111111111;
20'b00110100010101001110: color_data = 12'b111111111111;
20'b00110100010101001111: color_data = 12'b111111111111;
20'b00110100010101011000: color_data = 12'b111111111111;
20'b00110100010101011001: color_data = 12'b111111111111;
20'b00110100010101011010: color_data = 12'b111111111111;
20'b00110100010101011011: color_data = 12'b111111111111;
20'b00110100010101011100: color_data = 12'b111111111111;
20'b00110100010101011101: color_data = 12'b111111111111;
20'b00110100010101011110: color_data = 12'b111111111111;
20'b00110100010101011111: color_data = 12'b111111111111;
20'b00110100010101100000: color_data = 12'b111111111111;
20'b00110100010101100001: color_data = 12'b111111111111;
20'b00110100010101100010: color_data = 12'b111111111111;
20'b00110100010101100011: color_data = 12'b111111111111;
20'b00110100010101100100: color_data = 12'b111111111111;
20'b00110100010101100101: color_data = 12'b111111111111;
20'b00110100010101100110: color_data = 12'b111111111111;
20'b00110100010101100111: color_data = 12'b111111111111;
20'b00110100010101101100: color_data = 12'b111111111111;
20'b00110100010101101101: color_data = 12'b111111111111;
20'b00110100010101101110: color_data = 12'b111111111111;
20'b00110100010101101111: color_data = 12'b111111111111;
20'b00110100010101110000: color_data = 12'b111111111111;
20'b00110100010101110001: color_data = 12'b111111111111;
20'b00110100010101110010: color_data = 12'b111111111111;
20'b00110100010101110011: color_data = 12'b111111111111;
20'b00110100010101110100: color_data = 12'b111111111111;
20'b00110100010101110101: color_data = 12'b111111111111;
20'b00110100010101110110: color_data = 12'b111111111111;
20'b00110100010101110111: color_data = 12'b111111111111;
20'b00110100010101111000: color_data = 12'b111111111111;
20'b00110100010101111001: color_data = 12'b111111111111;
20'b00110100010101111010: color_data = 12'b111111111111;
20'b00110100010101111011: color_data = 12'b111111111111;
20'b00110100010110000100: color_data = 12'b111111111111;
20'b00110100010110000101: color_data = 12'b111111111111;
20'b00110100010110000110: color_data = 12'b111111111111;
20'b00110100010110000111: color_data = 12'b111111111111;
20'b00111000100100001000: color_data = 12'b111111111111;
20'b00111000100100001001: color_data = 12'b111111111111;
20'b00111000100100001010: color_data = 12'b111111111111;
20'b00111000100100001011: color_data = 12'b111111111111;
20'b00111000100100001100: color_data = 12'b111111111111;
20'b00111000100100100010: color_data = 12'b111111111111;
20'b00111000100100100011: color_data = 12'b111111111111;
20'b00111000100100100100: color_data = 12'b111111111111;
20'b00111000100100100101: color_data = 12'b111111111111;
20'b00111000100100100110: color_data = 12'b111111111111;
20'b00111000100100100111: color_data = 12'b111111111111;
20'b00111000100100101000: color_data = 12'b111111111111;
20'b00111000100100101001: color_data = 12'b111111111111;
20'b00111000100100101010: color_data = 12'b111111111111;
20'b00111000100100101011: color_data = 12'b111111111111;
20'b00111000100100101100: color_data = 12'b111111111111;
20'b00111000100100101101: color_data = 12'b111111111111;
20'b00111000100100101110: color_data = 12'b111111111111;
20'b00111000100100101111: color_data = 12'b111111111111;
20'b00111000100100110000: color_data = 12'b111111111111;
20'b00111000100100110001: color_data = 12'b111111111111;
20'b00111000100100110010: color_data = 12'b111111111111;
20'b00111000100100110011: color_data = 12'b111111111111;
20'b00111000100100110100: color_data = 12'b111111111111;
20'b00111000100100110101: color_data = 12'b111111111111;
20'b00111000100100111100: color_data = 12'b111111111111;
20'b00111000100100111101: color_data = 12'b111111111111;
20'b00111000100100111110: color_data = 12'b111111111111;
20'b00111000100100111111: color_data = 12'b111111111111;
20'b00111000100101000000: color_data = 12'b111111111111;
20'b00111000100101001011: color_data = 12'b111111111111;
20'b00111000100101001100: color_data = 12'b111111111111;
20'b00111000100101001101: color_data = 12'b111111111111;
20'b00111000100101001110: color_data = 12'b111111111111;
20'b00111000100101001111: color_data = 12'b111111111111;
20'b00111000100101010101: color_data = 12'b111111111111;
20'b00111000100101010110: color_data = 12'b111111111111;
20'b00111000100101010111: color_data = 12'b111111111111;
20'b00111000100101011000: color_data = 12'b111111111111;
20'b00111000100101011001: color_data = 12'b111111111111;
20'b00111000100101011010: color_data = 12'b111111111111;
20'b00111000100101011011: color_data = 12'b111111111111;
20'b00111000100101011100: color_data = 12'b111111111111;
20'b00111000100101011101: color_data = 12'b111111111111;
20'b00111000100101011110: color_data = 12'b111111111111;
20'b00111000100101011111: color_data = 12'b111111111111;
20'b00111000100101100000: color_data = 12'b111111111111;
20'b00111000100101100001: color_data = 12'b111111111111;
20'b00111000100101100010: color_data = 12'b111111111111;
20'b00111000100101100011: color_data = 12'b111111111111;
20'b00111000100101100100: color_data = 12'b111111111111;
20'b00111000100101100101: color_data = 12'b111111111111;
20'b00111000100101100110: color_data = 12'b111111111111;
20'b00111000100101100111: color_data = 12'b111111111111;
20'b00111000100101101000: color_data = 12'b111111111111;
20'b00111000100101101001: color_data = 12'b111111111111;
20'b00111000100101101111: color_data = 12'b111111111111;
20'b00111000100101110000: color_data = 12'b111111111111;
20'b00111000100101110001: color_data = 12'b111111111111;
20'b00111000100101110010: color_data = 12'b111111111111;
20'b00111000100101110011: color_data = 12'b111111111111;
20'b00111000100110001101: color_data = 12'b111111111111;
20'b00111000100110001110: color_data = 12'b111111111111;
20'b00111000100110001111: color_data = 12'b111111111111;
20'b00111000100110010000: color_data = 12'b111111111111;
20'b00111000100110010001: color_data = 12'b111111111111;
20'b00111000100110010010: color_data = 12'b111111111111;
20'b00111000100110010011: color_data = 12'b111111111111;
20'b00111000100110010100: color_data = 12'b111111111111;
20'b00111000100110010101: color_data = 12'b111111111111;
20'b00111000100110010110: color_data = 12'b111111111111;
20'b00111000100110010111: color_data = 12'b111111111111;
20'b00111000100110011000: color_data = 12'b111111111111;
20'b00111000100110011001: color_data = 12'b111111111111;
20'b00111000100110011010: color_data = 12'b111111111111;
20'b00111000100110011011: color_data = 12'b111111111111;
20'b00111000100110011100: color_data = 12'b111111111111;
20'b00111000100110011101: color_data = 12'b111111111111;
20'b00111000100110011110: color_data = 12'b111111111111;
20'b00111000100110011111: color_data = 12'b111111111111;
20'b00111000100110100000: color_data = 12'b111111111111;
20'b00111000110100001000: color_data = 12'b111111111111;
20'b00111000110100001001: color_data = 12'b111111111111;
20'b00111000110100001010: color_data = 12'b111111111111;
20'b00111000110100001011: color_data = 12'b111111111111;
20'b00111000110100001100: color_data = 12'b111111111111;
20'b00111000110100100010: color_data = 12'b111111111111;
20'b00111000110100100011: color_data = 12'b111111111111;
20'b00111000110100100100: color_data = 12'b111111111111;
20'b00111000110100100101: color_data = 12'b111111111111;
20'b00111000110100100110: color_data = 12'b111111111111;
20'b00111000110100100111: color_data = 12'b111111111111;
20'b00111000110100101000: color_data = 12'b111111111111;
20'b00111000110100101001: color_data = 12'b111111111111;
20'b00111000110100101010: color_data = 12'b111111111111;
20'b00111000110100101011: color_data = 12'b111111111111;
20'b00111000110100101100: color_data = 12'b111111111111;
20'b00111000110100101101: color_data = 12'b111111111111;
20'b00111000110100101110: color_data = 12'b111111111111;
20'b00111000110100101111: color_data = 12'b111111111111;
20'b00111000110100110000: color_data = 12'b111111111111;
20'b00111000110100110001: color_data = 12'b111111111111;
20'b00111000110100110010: color_data = 12'b111111111111;
20'b00111000110100110011: color_data = 12'b111111111111;
20'b00111000110100110100: color_data = 12'b111111111111;
20'b00111000110100110101: color_data = 12'b111111111111;
20'b00111000110100111100: color_data = 12'b111111111111;
20'b00111000110100111101: color_data = 12'b111111111111;
20'b00111000110100111110: color_data = 12'b111111111111;
20'b00111000110100111111: color_data = 12'b111111111111;
20'b00111000110101000000: color_data = 12'b111111111111;
20'b00111000110101001011: color_data = 12'b111111111111;
20'b00111000110101001100: color_data = 12'b111111111111;
20'b00111000110101001101: color_data = 12'b111111111111;
20'b00111000110101001110: color_data = 12'b111111111111;
20'b00111000110101001111: color_data = 12'b111111111111;
20'b00111000110101010101: color_data = 12'b111111111111;
20'b00111000110101010110: color_data = 12'b111111111111;
20'b00111000110101010111: color_data = 12'b111111111111;
20'b00111000110101011000: color_data = 12'b111111111111;
20'b00111000110101011001: color_data = 12'b111111111111;
20'b00111000110101011010: color_data = 12'b111111111111;
20'b00111000110101011011: color_data = 12'b111111111111;
20'b00111000110101011100: color_data = 12'b111111111111;
20'b00111000110101011101: color_data = 12'b111111111111;
20'b00111000110101011110: color_data = 12'b111111111111;
20'b00111000110101011111: color_data = 12'b111111111111;
20'b00111000110101100000: color_data = 12'b111111111111;
20'b00111000110101100001: color_data = 12'b111111111111;
20'b00111000110101100010: color_data = 12'b111111111111;
20'b00111000110101100011: color_data = 12'b111111111111;
20'b00111000110101100100: color_data = 12'b111111111111;
20'b00111000110101100101: color_data = 12'b111111111111;
20'b00111000110101100110: color_data = 12'b111111111111;
20'b00111000110101100111: color_data = 12'b111111111111;
20'b00111000110101101000: color_data = 12'b111111111111;
20'b00111000110101101001: color_data = 12'b111111111111;
20'b00111000110101101111: color_data = 12'b111111111111;
20'b00111000110101110000: color_data = 12'b111111111111;
20'b00111000110101110001: color_data = 12'b111111111111;
20'b00111000110101110010: color_data = 12'b111111111111;
20'b00111000110101110011: color_data = 12'b111111111111;
20'b00111000110110001101: color_data = 12'b111111111111;
20'b00111000110110001110: color_data = 12'b111111111111;
20'b00111000110110001111: color_data = 12'b111111111111;
20'b00111000110110010000: color_data = 12'b111111111111;
20'b00111000110110010001: color_data = 12'b111111111111;
20'b00111000110110010010: color_data = 12'b111111111111;
20'b00111000110110010011: color_data = 12'b111111111111;
20'b00111000110110010100: color_data = 12'b111111111111;
20'b00111000110110010101: color_data = 12'b111111111111;
20'b00111000110110010110: color_data = 12'b111111111111;
20'b00111000110110010111: color_data = 12'b111111111111;
20'b00111000110110011000: color_data = 12'b111111111111;
20'b00111000110110011001: color_data = 12'b111111111111;
20'b00111000110110011010: color_data = 12'b111111111111;
20'b00111000110110011011: color_data = 12'b111111111111;
20'b00111000110110011100: color_data = 12'b111111111111;
20'b00111000110110011101: color_data = 12'b111111111111;
20'b00111000110110011110: color_data = 12'b111111111111;
20'b00111000110110011111: color_data = 12'b111111111111;
20'b00111000110110100000: color_data = 12'b111111111111;
20'b00111001000100001000: color_data = 12'b111111111111;
20'b00111001000100001001: color_data = 12'b111111111111;
20'b00111001000100001010: color_data = 12'b111111111111;
20'b00111001000100001011: color_data = 12'b111111111111;
20'b00111001000100001100: color_data = 12'b111111111111;
20'b00111001000100100010: color_data = 12'b111111111111;
20'b00111001000100100011: color_data = 12'b111111111111;
20'b00111001000100100100: color_data = 12'b111111111111;
20'b00111001000100100101: color_data = 12'b111111111111;
20'b00111001000100100110: color_data = 12'b111111111111;
20'b00111001000100100111: color_data = 12'b111111111111;
20'b00111001000100101000: color_data = 12'b111111111111;
20'b00111001000100101001: color_data = 12'b111111111111;
20'b00111001000100101010: color_data = 12'b111111111111;
20'b00111001000100101011: color_data = 12'b111111111111;
20'b00111001000100101100: color_data = 12'b111111111111;
20'b00111001000100101101: color_data = 12'b111111111111;
20'b00111001000100101110: color_data = 12'b111111111111;
20'b00111001000100101111: color_data = 12'b111111111111;
20'b00111001000100110000: color_data = 12'b111111111111;
20'b00111001000100110001: color_data = 12'b111111111111;
20'b00111001000100110010: color_data = 12'b111111111111;
20'b00111001000100110011: color_data = 12'b111111111111;
20'b00111001000100110100: color_data = 12'b111111111111;
20'b00111001000100110101: color_data = 12'b111111111111;
20'b00111001000100111100: color_data = 12'b111111111111;
20'b00111001000100111101: color_data = 12'b111111111111;
20'b00111001000100111110: color_data = 12'b111111111111;
20'b00111001000100111111: color_data = 12'b111111111111;
20'b00111001000101000000: color_data = 12'b111111111111;
20'b00111001000101001011: color_data = 12'b111111111111;
20'b00111001000101001100: color_data = 12'b111111111111;
20'b00111001000101001101: color_data = 12'b111111111111;
20'b00111001000101001110: color_data = 12'b111111111111;
20'b00111001000101001111: color_data = 12'b111111111111;
20'b00111001000101010101: color_data = 12'b111111111111;
20'b00111001000101010110: color_data = 12'b111111111111;
20'b00111001000101010111: color_data = 12'b111111111111;
20'b00111001000101011000: color_data = 12'b111111111111;
20'b00111001000101011001: color_data = 12'b111111111111;
20'b00111001000101011010: color_data = 12'b111111111111;
20'b00111001000101011011: color_data = 12'b111111111111;
20'b00111001000101011100: color_data = 12'b111111111111;
20'b00111001000101011101: color_data = 12'b111111111111;
20'b00111001000101011110: color_data = 12'b111111111111;
20'b00111001000101011111: color_data = 12'b111111111111;
20'b00111001000101100000: color_data = 12'b111111111111;
20'b00111001000101100001: color_data = 12'b111111111111;
20'b00111001000101100010: color_data = 12'b111111111111;
20'b00111001000101100011: color_data = 12'b111111111111;
20'b00111001000101100100: color_data = 12'b111111111111;
20'b00111001000101100101: color_data = 12'b111111111111;
20'b00111001000101100110: color_data = 12'b111111111111;
20'b00111001000101100111: color_data = 12'b111111111111;
20'b00111001000101101000: color_data = 12'b111111111111;
20'b00111001000101101001: color_data = 12'b111111111111;
20'b00111001000101101111: color_data = 12'b111111111111;
20'b00111001000101110000: color_data = 12'b111111111111;
20'b00111001000101110001: color_data = 12'b111111111111;
20'b00111001000101110010: color_data = 12'b111111111111;
20'b00111001000101110011: color_data = 12'b111111111111;
20'b00111001000110001101: color_data = 12'b111111111111;
20'b00111001000110001110: color_data = 12'b111111111111;
20'b00111001000110001111: color_data = 12'b111111111111;
20'b00111001000110010000: color_data = 12'b111111111111;
20'b00111001000110010001: color_data = 12'b111111111111;
20'b00111001000110010010: color_data = 12'b111111111111;
20'b00111001000110010011: color_data = 12'b111111111111;
20'b00111001000110010100: color_data = 12'b111111111111;
20'b00111001000110010101: color_data = 12'b111111111111;
20'b00111001000110010110: color_data = 12'b111111111111;
20'b00111001000110010111: color_data = 12'b111111111111;
20'b00111001000110011000: color_data = 12'b111111111111;
20'b00111001000110011001: color_data = 12'b111111111111;
20'b00111001000110011010: color_data = 12'b111111111111;
20'b00111001000110011011: color_data = 12'b111111111111;
20'b00111001000110011100: color_data = 12'b111111111111;
20'b00111001000110011101: color_data = 12'b111111111111;
20'b00111001000110011110: color_data = 12'b111111111111;
20'b00111001000110011111: color_data = 12'b111111111111;
20'b00111001000110100000: color_data = 12'b111111111111;
20'b00111001010100001000: color_data = 12'b111111111111;
20'b00111001010100001001: color_data = 12'b111111111111;
20'b00111001010100001010: color_data = 12'b111111111111;
20'b00111001010100001011: color_data = 12'b111111111111;
20'b00111001010100001100: color_data = 12'b111111111111;
20'b00111001010100100010: color_data = 12'b111111111111;
20'b00111001010100100011: color_data = 12'b111111111111;
20'b00111001010100100100: color_data = 12'b111111111111;
20'b00111001010100100101: color_data = 12'b111111111111;
20'b00111001010100100110: color_data = 12'b111111111111;
20'b00111001010100100111: color_data = 12'b111111111111;
20'b00111001010100101000: color_data = 12'b111111111111;
20'b00111001010100101001: color_data = 12'b111111111111;
20'b00111001010100101010: color_data = 12'b111111111111;
20'b00111001010100101011: color_data = 12'b111111111111;
20'b00111001010100101100: color_data = 12'b111111111111;
20'b00111001010100101101: color_data = 12'b111111111111;
20'b00111001010100101110: color_data = 12'b111111111111;
20'b00111001010100101111: color_data = 12'b111111111111;
20'b00111001010100110000: color_data = 12'b111111111111;
20'b00111001010100110001: color_data = 12'b111111111111;
20'b00111001010100110010: color_data = 12'b111111111111;
20'b00111001010100110011: color_data = 12'b111111111111;
20'b00111001010100110100: color_data = 12'b111111111111;
20'b00111001010100110101: color_data = 12'b111111111111;
20'b00111001010100111100: color_data = 12'b111111111111;
20'b00111001010100111101: color_data = 12'b111111111111;
20'b00111001010100111110: color_data = 12'b111111111111;
20'b00111001010100111111: color_data = 12'b111111111111;
20'b00111001010101000000: color_data = 12'b111111111111;
20'b00111001010101001011: color_data = 12'b111111111111;
20'b00111001010101001100: color_data = 12'b111111111111;
20'b00111001010101001101: color_data = 12'b111111111111;
20'b00111001010101001110: color_data = 12'b111111111111;
20'b00111001010101001111: color_data = 12'b111111111111;
20'b00111001010101010101: color_data = 12'b111111111111;
20'b00111001010101010110: color_data = 12'b111111111111;
20'b00111001010101010111: color_data = 12'b111111111111;
20'b00111001010101011000: color_data = 12'b111111111111;
20'b00111001010101011001: color_data = 12'b111111111111;
20'b00111001010101011010: color_data = 12'b111111111111;
20'b00111001010101011011: color_data = 12'b111111111111;
20'b00111001010101011100: color_data = 12'b111111111111;
20'b00111001010101011101: color_data = 12'b111111111111;
20'b00111001010101011110: color_data = 12'b111111111111;
20'b00111001010101011111: color_data = 12'b111111111111;
20'b00111001010101100000: color_data = 12'b111111111111;
20'b00111001010101100001: color_data = 12'b111111111111;
20'b00111001010101100010: color_data = 12'b111111111111;
20'b00111001010101100011: color_data = 12'b111111111111;
20'b00111001010101100100: color_data = 12'b111111111111;
20'b00111001010101100101: color_data = 12'b111111111111;
20'b00111001010101100110: color_data = 12'b111111111111;
20'b00111001010101100111: color_data = 12'b111111111111;
20'b00111001010101101000: color_data = 12'b111111111111;
20'b00111001010101101001: color_data = 12'b111111111111;
20'b00111001010101101111: color_data = 12'b111111111111;
20'b00111001010101110000: color_data = 12'b111111111111;
20'b00111001010101110001: color_data = 12'b111111111111;
20'b00111001010101110010: color_data = 12'b111111111111;
20'b00111001010101110011: color_data = 12'b111111111111;
20'b00111001010110001101: color_data = 12'b111111111111;
20'b00111001010110001110: color_data = 12'b111111111111;
20'b00111001010110001111: color_data = 12'b111111111111;
20'b00111001010110010000: color_data = 12'b111111111111;
20'b00111001010110010001: color_data = 12'b111111111111;
20'b00111001010110010010: color_data = 12'b111111111111;
20'b00111001010110010011: color_data = 12'b111111111111;
20'b00111001010110010100: color_data = 12'b111111111111;
20'b00111001010110010101: color_data = 12'b111111111111;
20'b00111001010110010110: color_data = 12'b111111111111;
20'b00111001010110010111: color_data = 12'b111111111111;
20'b00111001010110011000: color_data = 12'b111111111111;
20'b00111001010110011001: color_data = 12'b111111111111;
20'b00111001010110011010: color_data = 12'b111111111111;
20'b00111001010110011011: color_data = 12'b111111111111;
20'b00111001010110011100: color_data = 12'b111111111111;
20'b00111001010110011101: color_data = 12'b111111111111;
20'b00111001010110011110: color_data = 12'b111111111111;
20'b00111001010110011111: color_data = 12'b111111111111;
20'b00111001010110100000: color_data = 12'b111111111111;
20'b00111001100100001000: color_data = 12'b111111111111;
20'b00111001100100001001: color_data = 12'b111111111111;
20'b00111001100100001010: color_data = 12'b111111111111;
20'b00111001100100001011: color_data = 12'b111111111111;
20'b00111001100100001100: color_data = 12'b111111111111;
20'b00111001100100100010: color_data = 12'b111111111111;
20'b00111001100100100011: color_data = 12'b111111111111;
20'b00111001100100100100: color_data = 12'b111111111111;
20'b00111001100100100101: color_data = 12'b111111111111;
20'b00111001100100100110: color_data = 12'b111111111111;
20'b00111001100100111100: color_data = 12'b111111111111;
20'b00111001100100111101: color_data = 12'b111111111111;
20'b00111001100100111110: color_data = 12'b111111111111;
20'b00111001100100111111: color_data = 12'b111111111111;
20'b00111001100101000000: color_data = 12'b111111111111;
20'b00111001100101001011: color_data = 12'b111111111111;
20'b00111001100101001100: color_data = 12'b111111111111;
20'b00111001100101001101: color_data = 12'b111111111111;
20'b00111001100101001110: color_data = 12'b111111111111;
20'b00111001100101001111: color_data = 12'b111111111111;
20'b00111001100101010101: color_data = 12'b111111111111;
20'b00111001100101010110: color_data = 12'b111111111111;
20'b00111001100101010111: color_data = 12'b111111111111;
20'b00111001100101011000: color_data = 12'b111111111111;
20'b00111001100101011001: color_data = 12'b111111111111;
20'b00111001100101101111: color_data = 12'b111111111111;
20'b00111001100101110000: color_data = 12'b111111111111;
20'b00111001100101110001: color_data = 12'b111111111111;
20'b00111001100101110010: color_data = 12'b111111111111;
20'b00111001100101110011: color_data = 12'b111111111111;
20'b00111001100110011101: color_data = 12'b111111111111;
20'b00111001100110011110: color_data = 12'b111111111111;
20'b00111001100110011111: color_data = 12'b111111111111;
20'b00111001100110100000: color_data = 12'b111111111111;
20'b00111001110100001000: color_data = 12'b111111111111;
20'b00111001110100001001: color_data = 12'b111111111111;
20'b00111001110100001010: color_data = 12'b111111111111;
20'b00111001110100001011: color_data = 12'b111111111111;
20'b00111001110100001100: color_data = 12'b111111111111;
20'b00111001110100100010: color_data = 12'b111111111111;
20'b00111001110100100011: color_data = 12'b111111111111;
20'b00111001110100100100: color_data = 12'b111111111111;
20'b00111001110100100101: color_data = 12'b111111111111;
20'b00111001110100100110: color_data = 12'b111111111111;
20'b00111001110100111100: color_data = 12'b111111111111;
20'b00111001110100111101: color_data = 12'b111111111111;
20'b00111001110100111110: color_data = 12'b111111111111;
20'b00111001110100111111: color_data = 12'b111111111111;
20'b00111001110101000000: color_data = 12'b111111111111;
20'b00111001110101001011: color_data = 12'b111111111111;
20'b00111001110101001100: color_data = 12'b111111111111;
20'b00111001110101001101: color_data = 12'b111111111111;
20'b00111001110101001110: color_data = 12'b111111111111;
20'b00111001110101001111: color_data = 12'b111111111111;
20'b00111001110101010101: color_data = 12'b111111111111;
20'b00111001110101010110: color_data = 12'b111111111111;
20'b00111001110101010111: color_data = 12'b111111111111;
20'b00111001110101011000: color_data = 12'b111111111111;
20'b00111001110101011001: color_data = 12'b111111111111;
20'b00111001110101101111: color_data = 12'b111111111111;
20'b00111001110101110000: color_data = 12'b111111111111;
20'b00111001110101110001: color_data = 12'b111111111111;
20'b00111001110101110010: color_data = 12'b111111111111;
20'b00111001110101110011: color_data = 12'b111111111111;
20'b00111001110110011101: color_data = 12'b111111111111;
20'b00111001110110011110: color_data = 12'b111111111111;
20'b00111001110110011111: color_data = 12'b111111111111;
20'b00111001110110100000: color_data = 12'b111111111111;
20'b00111010000100001000: color_data = 12'b111111111111;
20'b00111010000100001001: color_data = 12'b111111111111;
20'b00111010000100001010: color_data = 12'b111111111111;
20'b00111010000100001011: color_data = 12'b111111111111;
20'b00111010000100001100: color_data = 12'b111111111111;
20'b00111010000100100010: color_data = 12'b111111111111;
20'b00111010000100100011: color_data = 12'b111111111111;
20'b00111010000100100100: color_data = 12'b111111111111;
20'b00111010000100100101: color_data = 12'b111111111111;
20'b00111010000100100110: color_data = 12'b111111111111;
20'b00111010000100111100: color_data = 12'b111111111111;
20'b00111010000100111101: color_data = 12'b111111111111;
20'b00111010000100111110: color_data = 12'b111111111111;
20'b00111010000100111111: color_data = 12'b111111111111;
20'b00111010000101000000: color_data = 12'b111111111111;
20'b00111010000101001011: color_data = 12'b111111111111;
20'b00111010000101001100: color_data = 12'b111111111111;
20'b00111010000101001101: color_data = 12'b111111111111;
20'b00111010000101001110: color_data = 12'b111111111111;
20'b00111010000101001111: color_data = 12'b111111111111;
20'b00111010000101010101: color_data = 12'b111111111111;
20'b00111010000101010110: color_data = 12'b111111111111;
20'b00111010000101010111: color_data = 12'b111111111111;
20'b00111010000101011000: color_data = 12'b111111111111;
20'b00111010000101011001: color_data = 12'b111111111111;
20'b00111010000101101111: color_data = 12'b111111111111;
20'b00111010000101110000: color_data = 12'b111111111111;
20'b00111010000101110001: color_data = 12'b111111111111;
20'b00111010000101110010: color_data = 12'b111111111111;
20'b00111010000101110011: color_data = 12'b111111111111;
20'b00111010000110011101: color_data = 12'b111111111111;
20'b00111010000110011110: color_data = 12'b111111111111;
20'b00111010000110011111: color_data = 12'b111111111111;
20'b00111010000110100000: color_data = 12'b111111111111;
20'b00111010010011111011: color_data = 12'b111111111111;
20'b00111010010011111100: color_data = 12'b111111111111;
20'b00111010010011111101: color_data = 12'b111111111111;
20'b00111010010011111110: color_data = 12'b111111111111;
20'b00111010010011111111: color_data = 12'b111111111111;
20'b00111010010100000000: color_data = 12'b111111111111;
20'b00111010010100000001: color_data = 12'b111111111111;
20'b00111010010100001000: color_data = 12'b111111111111;
20'b00111010010100001001: color_data = 12'b111111111111;
20'b00111010010100001010: color_data = 12'b111111111111;
20'b00111010010100001011: color_data = 12'b111111111111;
20'b00111010010100001100: color_data = 12'b111111111111;
20'b00111010010100100010: color_data = 12'b111111111111;
20'b00111010010100100011: color_data = 12'b111111111111;
20'b00111010010100100100: color_data = 12'b111111111111;
20'b00111010010100100101: color_data = 12'b111111111111;
20'b00111010010100100110: color_data = 12'b111111111111;
20'b00111010010100111100: color_data = 12'b111111111111;
20'b00111010010100111101: color_data = 12'b111111111111;
20'b00111010010100111110: color_data = 12'b111111111111;
20'b00111010010100111111: color_data = 12'b111111111111;
20'b00111010010101000000: color_data = 12'b111111111111;
20'b00111010010101001011: color_data = 12'b111111111111;
20'b00111010010101001100: color_data = 12'b111111111111;
20'b00111010010101001101: color_data = 12'b111111111111;
20'b00111010010101001110: color_data = 12'b111111111111;
20'b00111010010101001111: color_data = 12'b111111111111;
20'b00111010010101010101: color_data = 12'b111111111111;
20'b00111010010101010110: color_data = 12'b111111111111;
20'b00111010010101010111: color_data = 12'b111111111111;
20'b00111010010101011000: color_data = 12'b111111111111;
20'b00111010010101011001: color_data = 12'b111111111111;
20'b00111010010101101111: color_data = 12'b111111111111;
20'b00111010010101110000: color_data = 12'b111111111111;
20'b00111010010101110001: color_data = 12'b111111111111;
20'b00111010010101110010: color_data = 12'b111111111111;
20'b00111010010101110011: color_data = 12'b111111111111;
20'b00111010010110011101: color_data = 12'b111111111111;
20'b00111010010110011110: color_data = 12'b111111111111;
20'b00111010010110011111: color_data = 12'b111111111111;
20'b00111010010110100000: color_data = 12'b111111111111;
20'b00111010100011111011: color_data = 12'b111111111111;
20'b00111010100011111100: color_data = 12'b111111111111;
20'b00111010100011111101: color_data = 12'b111111111111;
20'b00111010100011111110: color_data = 12'b111111111111;
20'b00111010100011111111: color_data = 12'b111111111111;
20'b00111010100100000000: color_data = 12'b111111111111;
20'b00111010100100000001: color_data = 12'b111111111111;
20'b00111010100100001000: color_data = 12'b111111111111;
20'b00111010100100001001: color_data = 12'b111111111111;
20'b00111010100100001010: color_data = 12'b111111111111;
20'b00111010100100001011: color_data = 12'b111111111111;
20'b00111010100100001100: color_data = 12'b111111111111;
20'b00111010100100100010: color_data = 12'b111111111111;
20'b00111010100100100011: color_data = 12'b111111111111;
20'b00111010100100100100: color_data = 12'b111111111111;
20'b00111010100100100101: color_data = 12'b111111111111;
20'b00111010100100100110: color_data = 12'b111111111111;
20'b00111010100100100111: color_data = 12'b111111111111;
20'b00111010100100101000: color_data = 12'b111111111111;
20'b00111010100100101001: color_data = 12'b111111111111;
20'b00111010100100101010: color_data = 12'b111111111111;
20'b00111010100100101011: color_data = 12'b111111111111;
20'b00111010100100101100: color_data = 12'b111111111111;
20'b00111010100100101101: color_data = 12'b111111111111;
20'b00111010100100101110: color_data = 12'b111111111111;
20'b00111010100100101111: color_data = 12'b111111111111;
20'b00111010100100110000: color_data = 12'b111111111111;
20'b00111010100100110001: color_data = 12'b111111111111;
20'b00111010100100110010: color_data = 12'b111111111111;
20'b00111010100100110011: color_data = 12'b111111111111;
20'b00111010100100110100: color_data = 12'b111111111111;
20'b00111010100100110101: color_data = 12'b111111111111;
20'b00111010100100111100: color_data = 12'b111111111111;
20'b00111010100100111101: color_data = 12'b111111111111;
20'b00111010100100111110: color_data = 12'b111111111111;
20'b00111010100100111111: color_data = 12'b111111111111;
20'b00111010100101000000: color_data = 12'b111111111111;
20'b00111010100101001011: color_data = 12'b111111111111;
20'b00111010100101001100: color_data = 12'b111111111111;
20'b00111010100101001101: color_data = 12'b111111111111;
20'b00111010100101001110: color_data = 12'b111111111111;
20'b00111010100101001111: color_data = 12'b111111111111;
20'b00111010100101010101: color_data = 12'b111111111111;
20'b00111010100101010110: color_data = 12'b111111111111;
20'b00111010100101010111: color_data = 12'b111111111111;
20'b00111010100101011000: color_data = 12'b111111111111;
20'b00111010100101011001: color_data = 12'b111111111111;
20'b00111010100101011010: color_data = 12'b111111111111;
20'b00111010100101011011: color_data = 12'b111111111111;
20'b00111010100101011100: color_data = 12'b111111111111;
20'b00111010100101011101: color_data = 12'b111111111111;
20'b00111010100101011110: color_data = 12'b111111111111;
20'b00111010100101011111: color_data = 12'b111111111111;
20'b00111010100101100000: color_data = 12'b111111111111;
20'b00111010100101100001: color_data = 12'b111111111111;
20'b00111010100101100010: color_data = 12'b111111111111;
20'b00111010100101100011: color_data = 12'b111111111111;
20'b00111010100101100100: color_data = 12'b111111111111;
20'b00111010100101100101: color_data = 12'b111111111111;
20'b00111010100101100110: color_data = 12'b111111111111;
20'b00111010100101100111: color_data = 12'b111111111111;
20'b00111010100101101000: color_data = 12'b111111111111;
20'b00111010100101101001: color_data = 12'b111111111111;
20'b00111010100101101111: color_data = 12'b111111111111;
20'b00111010100101110000: color_data = 12'b111111111111;
20'b00111010100101110001: color_data = 12'b111111111111;
20'b00111010100101110010: color_data = 12'b111111111111;
20'b00111010100101110011: color_data = 12'b111111111111;
20'b00111010100110001101: color_data = 12'b111111111111;
20'b00111010100110001110: color_data = 12'b111111111111;
20'b00111010100110001111: color_data = 12'b111111111111;
20'b00111010100110010000: color_data = 12'b111111111111;
20'b00111010100110010001: color_data = 12'b111111111111;
20'b00111010100110010010: color_data = 12'b111111111111;
20'b00111010100110010011: color_data = 12'b111111111111;
20'b00111010100110010100: color_data = 12'b111111111111;
20'b00111010100110010101: color_data = 12'b111111111111;
20'b00111010100110010110: color_data = 12'b111111111111;
20'b00111010100110010111: color_data = 12'b111111111111;
20'b00111010100110011000: color_data = 12'b111111111111;
20'b00111010100110011001: color_data = 12'b111111111111;
20'b00111010100110011010: color_data = 12'b111111111111;
20'b00111010100110011011: color_data = 12'b111111111111;
20'b00111010100110011100: color_data = 12'b111111111111;
20'b00111010100110011101: color_data = 12'b111111111111;
20'b00111010100110011110: color_data = 12'b111111111111;
20'b00111010100110011111: color_data = 12'b111111111111;
20'b00111010100110100000: color_data = 12'b111111111111;
20'b00111010110011111011: color_data = 12'b111111111111;
20'b00111010110011111100: color_data = 12'b111111111111;
20'b00111010110011111101: color_data = 12'b111111111111;
20'b00111010110011111110: color_data = 12'b111111111111;
20'b00111010110011111111: color_data = 12'b111111111111;
20'b00111010110100000000: color_data = 12'b111111111111;
20'b00111010110100000001: color_data = 12'b111111111111;
20'b00111010110100001000: color_data = 12'b111111111111;
20'b00111010110100001001: color_data = 12'b111111111111;
20'b00111010110100001010: color_data = 12'b111111111111;
20'b00111010110100001011: color_data = 12'b111111111111;
20'b00111010110100001100: color_data = 12'b111111111111;
20'b00111010110100100010: color_data = 12'b111111111111;
20'b00111010110100100011: color_data = 12'b111111111111;
20'b00111010110100100100: color_data = 12'b111111111111;
20'b00111010110100100101: color_data = 12'b111111111111;
20'b00111010110100100110: color_data = 12'b111111111111;
20'b00111010110100100111: color_data = 12'b111111111111;
20'b00111010110100101000: color_data = 12'b111111111111;
20'b00111010110100101001: color_data = 12'b111111111111;
20'b00111010110100101010: color_data = 12'b111111111111;
20'b00111010110100101011: color_data = 12'b111111111111;
20'b00111010110100101100: color_data = 12'b111111111111;
20'b00111010110100101101: color_data = 12'b111111111111;
20'b00111010110100101110: color_data = 12'b111111111111;
20'b00111010110100101111: color_data = 12'b111111111111;
20'b00111010110100110000: color_data = 12'b111111111111;
20'b00111010110100110001: color_data = 12'b111111111111;
20'b00111010110100110010: color_data = 12'b111111111111;
20'b00111010110100110011: color_data = 12'b111111111111;
20'b00111010110100110100: color_data = 12'b111111111111;
20'b00111010110100110101: color_data = 12'b111111111111;
20'b00111010110100111100: color_data = 12'b111111111111;
20'b00111010110100111101: color_data = 12'b111111111111;
20'b00111010110100111110: color_data = 12'b111111111111;
20'b00111010110100111111: color_data = 12'b111111111111;
20'b00111010110101000000: color_data = 12'b111111111111;
20'b00111010110101001011: color_data = 12'b111111111111;
20'b00111010110101001100: color_data = 12'b111111111111;
20'b00111010110101001101: color_data = 12'b111111111111;
20'b00111010110101001110: color_data = 12'b111111111111;
20'b00111010110101001111: color_data = 12'b111111111111;
20'b00111010110101010101: color_data = 12'b111111111111;
20'b00111010110101010110: color_data = 12'b111111111111;
20'b00111010110101010111: color_data = 12'b111111111111;
20'b00111010110101011000: color_data = 12'b111111111111;
20'b00111010110101011001: color_data = 12'b111111111111;
20'b00111010110101011010: color_data = 12'b111111111111;
20'b00111010110101011011: color_data = 12'b111111111111;
20'b00111010110101011100: color_data = 12'b111111111111;
20'b00111010110101011101: color_data = 12'b111111111111;
20'b00111010110101011110: color_data = 12'b111111111111;
20'b00111010110101011111: color_data = 12'b111111111111;
20'b00111010110101100000: color_data = 12'b111111111111;
20'b00111010110101100001: color_data = 12'b111111111111;
20'b00111010110101100010: color_data = 12'b111111111111;
20'b00111010110101100011: color_data = 12'b111111111111;
20'b00111010110101100100: color_data = 12'b111111111111;
20'b00111010110101100101: color_data = 12'b111111111111;
20'b00111010110101100110: color_data = 12'b111111111111;
20'b00111010110101100111: color_data = 12'b111111111111;
20'b00111010110101101000: color_data = 12'b111111111111;
20'b00111010110101101001: color_data = 12'b111111111111;
20'b00111010110101101111: color_data = 12'b111111111111;
20'b00111010110101110000: color_data = 12'b111111111111;
20'b00111010110101110001: color_data = 12'b111111111111;
20'b00111010110101110010: color_data = 12'b111111111111;
20'b00111010110101110011: color_data = 12'b111111111111;
20'b00111010110110001101: color_data = 12'b111111111111;
20'b00111010110110001110: color_data = 12'b111111111111;
20'b00111010110110001111: color_data = 12'b111111111111;
20'b00111010110110010000: color_data = 12'b111111111111;
20'b00111010110110010001: color_data = 12'b111111111111;
20'b00111010110110010010: color_data = 12'b111111111111;
20'b00111010110110010011: color_data = 12'b111111111111;
20'b00111010110110010100: color_data = 12'b111111111111;
20'b00111010110110010101: color_data = 12'b111111111111;
20'b00111010110110010110: color_data = 12'b111111111111;
20'b00111010110110010111: color_data = 12'b111111111111;
20'b00111010110110011000: color_data = 12'b111111111111;
20'b00111010110110011001: color_data = 12'b111111111111;
20'b00111010110110011010: color_data = 12'b111111111111;
20'b00111010110110011011: color_data = 12'b111111111111;
20'b00111010110110011100: color_data = 12'b111111111111;
20'b00111010110110011101: color_data = 12'b111111111111;
20'b00111010110110011110: color_data = 12'b111111111111;
20'b00111010110110011111: color_data = 12'b111111111111;
20'b00111010110110100000: color_data = 12'b111111111111;
20'b00111011000011111011: color_data = 12'b111111111111;
20'b00111011000011111100: color_data = 12'b111111111111;
20'b00111011000011111101: color_data = 12'b111111111111;
20'b00111011000011111110: color_data = 12'b111111111111;
20'b00111011000011111111: color_data = 12'b111111111111;
20'b00111011000100000000: color_data = 12'b111111111111;
20'b00111011000100000001: color_data = 12'b111111111111;
20'b00111011000100001000: color_data = 12'b111111111111;
20'b00111011000100001001: color_data = 12'b111111111111;
20'b00111011000100001010: color_data = 12'b111111111111;
20'b00111011000100001011: color_data = 12'b111111111111;
20'b00111011000100001100: color_data = 12'b111111111111;
20'b00111011000100100010: color_data = 12'b111111111111;
20'b00111011000100100011: color_data = 12'b111111111111;
20'b00111011000100100100: color_data = 12'b111111111111;
20'b00111011000100100101: color_data = 12'b111111111111;
20'b00111011000100100110: color_data = 12'b111111111111;
20'b00111011000100100111: color_data = 12'b111111111111;
20'b00111011000100101000: color_data = 12'b111111111111;
20'b00111011000100101001: color_data = 12'b111111111111;
20'b00111011000100101010: color_data = 12'b111111111111;
20'b00111011000100101011: color_data = 12'b111111111111;
20'b00111011000100101100: color_data = 12'b111111111111;
20'b00111011000100101101: color_data = 12'b111111111111;
20'b00111011000100101110: color_data = 12'b111111111111;
20'b00111011000100101111: color_data = 12'b111111111111;
20'b00111011000100110000: color_data = 12'b111111111111;
20'b00111011000100110001: color_data = 12'b111111111111;
20'b00111011000100110010: color_data = 12'b111111111111;
20'b00111011000100110011: color_data = 12'b111111111111;
20'b00111011000100110100: color_data = 12'b111111111111;
20'b00111011000100110101: color_data = 12'b111111111111;
20'b00111011000100111100: color_data = 12'b111111111111;
20'b00111011000100111101: color_data = 12'b111111111111;
20'b00111011000100111110: color_data = 12'b111111111111;
20'b00111011000100111111: color_data = 12'b111111111111;
20'b00111011000101000000: color_data = 12'b111111111111;
20'b00111011000101001011: color_data = 12'b111111111111;
20'b00111011000101001100: color_data = 12'b111111111111;
20'b00111011000101001101: color_data = 12'b111111111111;
20'b00111011000101001110: color_data = 12'b111111111111;
20'b00111011000101001111: color_data = 12'b111111111111;
20'b00111011000101010101: color_data = 12'b111111111111;
20'b00111011000101010110: color_data = 12'b111111111111;
20'b00111011000101010111: color_data = 12'b111111111111;
20'b00111011000101011000: color_data = 12'b111111111111;
20'b00111011000101011001: color_data = 12'b111111111111;
20'b00111011000101011010: color_data = 12'b111111111111;
20'b00111011000101011011: color_data = 12'b111111111111;
20'b00111011000101011100: color_data = 12'b111111111111;
20'b00111011000101011101: color_data = 12'b111111111111;
20'b00111011000101011110: color_data = 12'b111111111111;
20'b00111011000101011111: color_data = 12'b111111111111;
20'b00111011000101100000: color_data = 12'b111111111111;
20'b00111011000101100001: color_data = 12'b111111111111;
20'b00111011000101100010: color_data = 12'b111111111111;
20'b00111011000101100011: color_data = 12'b111111111111;
20'b00111011000101100100: color_data = 12'b111111111111;
20'b00111011000101100101: color_data = 12'b111111111111;
20'b00111011000101100110: color_data = 12'b111111111111;
20'b00111011000101100111: color_data = 12'b111111111111;
20'b00111011000101101000: color_data = 12'b111111111111;
20'b00111011000101101001: color_data = 12'b111111111111;
20'b00111011000101101111: color_data = 12'b111111111111;
20'b00111011000101110000: color_data = 12'b111111111111;
20'b00111011000101110001: color_data = 12'b111111111111;
20'b00111011000101110010: color_data = 12'b111111111111;
20'b00111011000101110011: color_data = 12'b111111111111;
20'b00111011000110001101: color_data = 12'b111111111111;
20'b00111011000110001110: color_data = 12'b111111111111;
20'b00111011000110001111: color_data = 12'b111111111111;
20'b00111011000110010000: color_data = 12'b111111111111;
20'b00111011000110010001: color_data = 12'b111111111111;
20'b00111011000110010010: color_data = 12'b111111111111;
20'b00111011000110010011: color_data = 12'b111111111111;
20'b00111011000110010100: color_data = 12'b111111111111;
20'b00111011000110010101: color_data = 12'b111111111111;
20'b00111011000110010110: color_data = 12'b111111111111;
20'b00111011000110010111: color_data = 12'b111111111111;
20'b00111011000110011000: color_data = 12'b111111111111;
20'b00111011000110011001: color_data = 12'b111111111111;
20'b00111011000110011010: color_data = 12'b111111111111;
20'b00111011000110011011: color_data = 12'b111111111111;
20'b00111011000110011100: color_data = 12'b111111111111;
20'b00111011000110011101: color_data = 12'b111111111111;
20'b00111011000110011110: color_data = 12'b111111111111;
20'b00111011000110011111: color_data = 12'b111111111111;
20'b00111011000110100000: color_data = 12'b111111111111;
20'b00111011010011111011: color_data = 12'b111111111111;
20'b00111011010011111100: color_data = 12'b111111111111;
20'b00111011010011111101: color_data = 12'b111111111111;
20'b00111011010011111110: color_data = 12'b111111111111;
20'b00111011010011111111: color_data = 12'b111111111111;
20'b00111011010100000000: color_data = 12'b111111111111;
20'b00111011010100000001: color_data = 12'b111111111111;
20'b00111011010100001000: color_data = 12'b111111111111;
20'b00111011010100001001: color_data = 12'b111111111111;
20'b00111011010100001010: color_data = 12'b111111111111;
20'b00111011010100001011: color_data = 12'b111111111111;
20'b00111011010100001100: color_data = 12'b111111111111;
20'b00111011010100100010: color_data = 12'b111111111111;
20'b00111011010100100011: color_data = 12'b111111111111;
20'b00111011010100100100: color_data = 12'b111111111111;
20'b00111011010100100101: color_data = 12'b111111111111;
20'b00111011010100100110: color_data = 12'b111111111111;
20'b00111011010100100111: color_data = 12'b111111111111;
20'b00111011010100101000: color_data = 12'b111111111111;
20'b00111011010100101001: color_data = 12'b111111111111;
20'b00111011010100101010: color_data = 12'b111111111111;
20'b00111011010100101011: color_data = 12'b111111111111;
20'b00111011010100101100: color_data = 12'b111111111111;
20'b00111011010100101101: color_data = 12'b111111111111;
20'b00111011010100101110: color_data = 12'b111111111111;
20'b00111011010100101111: color_data = 12'b111111111111;
20'b00111011010100110000: color_data = 12'b111111111111;
20'b00111011010100110001: color_data = 12'b111111111111;
20'b00111011010100110010: color_data = 12'b111111111111;
20'b00111011010100110011: color_data = 12'b111111111111;
20'b00111011010100110100: color_data = 12'b111111111111;
20'b00111011010100110101: color_data = 12'b111111111111;
20'b00111011010100111100: color_data = 12'b111111111111;
20'b00111011010100111101: color_data = 12'b111111111111;
20'b00111011010100111110: color_data = 12'b111111111111;
20'b00111011010100111111: color_data = 12'b111111111111;
20'b00111011010101000000: color_data = 12'b111111111111;
20'b00111011010101001011: color_data = 12'b111111111111;
20'b00111011010101001100: color_data = 12'b111111111111;
20'b00111011010101001101: color_data = 12'b111111111111;
20'b00111011010101001110: color_data = 12'b111111111111;
20'b00111011010101001111: color_data = 12'b111111111111;
20'b00111011010101010101: color_data = 12'b111111111111;
20'b00111011010101010110: color_data = 12'b111111111111;
20'b00111011010101010111: color_data = 12'b111111111111;
20'b00111011010101011000: color_data = 12'b111111111111;
20'b00111011010101011001: color_data = 12'b111111111111;
20'b00111011010101011010: color_data = 12'b111111111111;
20'b00111011010101011011: color_data = 12'b111111111111;
20'b00111011010101011100: color_data = 12'b111111111111;
20'b00111011010101011101: color_data = 12'b111111111111;
20'b00111011010101011110: color_data = 12'b111111111111;
20'b00111011010101011111: color_data = 12'b111111111111;
20'b00111011010101100000: color_data = 12'b111111111111;
20'b00111011010101100001: color_data = 12'b111111111111;
20'b00111011010101100010: color_data = 12'b111111111111;
20'b00111011010101100011: color_data = 12'b111111111111;
20'b00111011010101100100: color_data = 12'b111111111111;
20'b00111011010101100101: color_data = 12'b111111111111;
20'b00111011010101100110: color_data = 12'b111111111111;
20'b00111011010101100111: color_data = 12'b111111111111;
20'b00111011010101101000: color_data = 12'b111111111111;
20'b00111011010101101001: color_data = 12'b111111111111;
20'b00111011010101101111: color_data = 12'b111111111111;
20'b00111011010101110000: color_data = 12'b111111111111;
20'b00111011010101110001: color_data = 12'b111111111111;
20'b00111011010101110010: color_data = 12'b111111111111;
20'b00111011010101110011: color_data = 12'b111111111111;
20'b00111011010110001101: color_data = 12'b111111111111;
20'b00111011010110001110: color_data = 12'b111111111111;
20'b00111011010110001111: color_data = 12'b111111111111;
20'b00111011010110010000: color_data = 12'b111111111111;
20'b00111011010110010001: color_data = 12'b111111111111;
20'b00111011010110010010: color_data = 12'b111111111111;
20'b00111011010110010011: color_data = 12'b111111111111;
20'b00111011010110010100: color_data = 12'b111111111111;
20'b00111011010110010101: color_data = 12'b111111111111;
20'b00111011010110010110: color_data = 12'b111111111111;
20'b00111011010110010111: color_data = 12'b111111111111;
20'b00111011010110011000: color_data = 12'b111111111111;
20'b00111011010110011001: color_data = 12'b111111111111;
20'b00111011010110011010: color_data = 12'b111111111111;
20'b00111011010110011011: color_data = 12'b111111111111;
20'b00111011010110011100: color_data = 12'b111111111111;
20'b00111011010110011101: color_data = 12'b111111111111;
20'b00111011010110011110: color_data = 12'b111111111111;
20'b00111011010110011111: color_data = 12'b111111111111;
20'b00111011010110100000: color_data = 12'b111111111111;
20'b00111011100011111011: color_data = 12'b111111111111;
20'b00111011100011111100: color_data = 12'b111111111111;
20'b00111011100011111101: color_data = 12'b111111111111;
20'b00111011100011111110: color_data = 12'b111111111111;
20'b00111011100011111111: color_data = 12'b111111111111;
20'b00111011100100000000: color_data = 12'b111111111111;
20'b00111011100100000001: color_data = 12'b111111111111;
20'b00111011100100001000: color_data = 12'b111111111111;
20'b00111011100100001001: color_data = 12'b111111111111;
20'b00111011100100001010: color_data = 12'b111111111111;
20'b00111011100100001011: color_data = 12'b111111111111;
20'b00111011100100001100: color_data = 12'b111111111111;
20'b00111011100100100010: color_data = 12'b111111111111;
20'b00111011100100100011: color_data = 12'b111111111111;
20'b00111011100100100100: color_data = 12'b111111111111;
20'b00111011100100100101: color_data = 12'b111111111111;
20'b00111011100100100110: color_data = 12'b111111111111;
20'b00111011100100100111: color_data = 12'b111111111111;
20'b00111011100100101000: color_data = 12'b111111111111;
20'b00111011100100101001: color_data = 12'b111111111111;
20'b00111011100100101010: color_data = 12'b111111111111;
20'b00111011100100101011: color_data = 12'b111111111111;
20'b00111011100100101100: color_data = 12'b111111111111;
20'b00111011100100101101: color_data = 12'b111111111111;
20'b00111011100100101110: color_data = 12'b111111111111;
20'b00111011100100101111: color_data = 12'b111111111111;
20'b00111011100100110000: color_data = 12'b111111111111;
20'b00111011100100110001: color_data = 12'b111111111111;
20'b00111011100100110010: color_data = 12'b111111111111;
20'b00111011100100110011: color_data = 12'b111111111111;
20'b00111011100100110100: color_data = 12'b111111111111;
20'b00111011100100110101: color_data = 12'b111111111111;
20'b00111011100100111100: color_data = 12'b111111111111;
20'b00111011100100111101: color_data = 12'b111111111111;
20'b00111011100100111110: color_data = 12'b111111111111;
20'b00111011100100111111: color_data = 12'b111111111111;
20'b00111011100101000000: color_data = 12'b111111111111;
20'b00111011100101001011: color_data = 12'b111111111111;
20'b00111011100101001100: color_data = 12'b111111111111;
20'b00111011100101001101: color_data = 12'b111111111111;
20'b00111011100101001110: color_data = 12'b111111111111;
20'b00111011100101001111: color_data = 12'b111111111111;
20'b00111011100101010101: color_data = 12'b111111111111;
20'b00111011100101010110: color_data = 12'b111111111111;
20'b00111011100101010111: color_data = 12'b111111111111;
20'b00111011100101011000: color_data = 12'b111111111111;
20'b00111011100101011001: color_data = 12'b111111111111;
20'b00111011100101011010: color_data = 12'b111111111111;
20'b00111011100101011011: color_data = 12'b111111111111;
20'b00111011100101011100: color_data = 12'b111111111111;
20'b00111011100101011101: color_data = 12'b111111111111;
20'b00111011100101011110: color_data = 12'b111111111111;
20'b00111011100101011111: color_data = 12'b111111111111;
20'b00111011100101100000: color_data = 12'b111111111111;
20'b00111011100101100001: color_data = 12'b111111111111;
20'b00111011100101100010: color_data = 12'b111111111111;
20'b00111011100101100011: color_data = 12'b111111111111;
20'b00111011100101100100: color_data = 12'b111111111111;
20'b00111011100101100101: color_data = 12'b111111111111;
20'b00111011100101100110: color_data = 12'b111111111111;
20'b00111011100101100111: color_data = 12'b111111111111;
20'b00111011100101101000: color_data = 12'b111111111111;
20'b00111011100101101001: color_data = 12'b111111111111;
20'b00111011100101101111: color_data = 12'b111111111111;
20'b00111011100101110000: color_data = 12'b111111111111;
20'b00111011100101110001: color_data = 12'b111111111111;
20'b00111011100101110010: color_data = 12'b111111111111;
20'b00111011100101110011: color_data = 12'b111111111111;
20'b00111011100110001101: color_data = 12'b111111111111;
20'b00111011100110001110: color_data = 12'b111111111111;
20'b00111011100110001111: color_data = 12'b111111111111;
20'b00111011100110010000: color_data = 12'b111111111111;
20'b00111011100110010001: color_data = 12'b111111111111;
20'b00111011100110010010: color_data = 12'b111111111111;
20'b00111011100110010011: color_data = 12'b111111111111;
20'b00111011100110010100: color_data = 12'b111111111111;
20'b00111011100110010101: color_data = 12'b111111111111;
20'b00111011100110010110: color_data = 12'b111111111111;
20'b00111011100110010111: color_data = 12'b111111111111;
20'b00111011100110011000: color_data = 12'b111111111111;
20'b00111011100110011001: color_data = 12'b111111111111;
20'b00111011100110011010: color_data = 12'b111111111111;
20'b00111011100110011011: color_data = 12'b111111111111;
20'b00111011100110011100: color_data = 12'b111111111111;
20'b00111011100110011101: color_data = 12'b111111111111;
20'b00111011100110011110: color_data = 12'b111111111111;
20'b00111011100110011111: color_data = 12'b111111111111;
20'b00111011100110100000: color_data = 12'b111111111111;
20'b00111011110011111011: color_data = 12'b111111111111;
20'b00111011110011111100: color_data = 12'b111111111111;
20'b00111011110011111101: color_data = 12'b111111111111;
20'b00111011110011111110: color_data = 12'b111111111111;
20'b00111011110011111111: color_data = 12'b111111111111;
20'b00111011110100000000: color_data = 12'b111111111111;
20'b00111011110100000001: color_data = 12'b111111111111;
20'b00111011110100001000: color_data = 12'b111111111111;
20'b00111011110100001001: color_data = 12'b111111111111;
20'b00111011110100001010: color_data = 12'b111111111111;
20'b00111011110100001011: color_data = 12'b111111111111;
20'b00111011110100001100: color_data = 12'b111111111111;
20'b00111011110100100010: color_data = 12'b111111111111;
20'b00111011110100100011: color_data = 12'b111111111111;
20'b00111011110100100100: color_data = 12'b111111111111;
20'b00111011110100100101: color_data = 12'b111111111111;
20'b00111011110100100110: color_data = 12'b111111111111;
20'b00111011110100100111: color_data = 12'b111111111111;
20'b00111011110100101000: color_data = 12'b111111111111;
20'b00111011110100101001: color_data = 12'b111111111111;
20'b00111011110100101010: color_data = 12'b111111111111;
20'b00111011110100101011: color_data = 12'b111111111111;
20'b00111011110100101100: color_data = 12'b111111111111;
20'b00111011110100101101: color_data = 12'b111111111111;
20'b00111011110100101110: color_data = 12'b111111111111;
20'b00111011110100101111: color_data = 12'b111111111111;
20'b00111011110100110000: color_data = 12'b111111111111;
20'b00111011110100110001: color_data = 12'b111111111111;
20'b00111011110100110010: color_data = 12'b111111111111;
20'b00111011110100110011: color_data = 12'b111111111111;
20'b00111011110100110100: color_data = 12'b111111111111;
20'b00111011110100110101: color_data = 12'b111111111111;
20'b00111011110100111100: color_data = 12'b111111111111;
20'b00111011110100111101: color_data = 12'b111111111111;
20'b00111011110100111110: color_data = 12'b111111111111;
20'b00111011110100111111: color_data = 12'b111111111111;
20'b00111011110101000000: color_data = 12'b111111111111;
20'b00111011110101001011: color_data = 12'b111111111111;
20'b00111011110101001100: color_data = 12'b111111111111;
20'b00111011110101001101: color_data = 12'b111111111111;
20'b00111011110101001110: color_data = 12'b111111111111;
20'b00111011110101001111: color_data = 12'b111111111111;
20'b00111011110101010101: color_data = 12'b111111111111;
20'b00111011110101010110: color_data = 12'b111111111111;
20'b00111011110101010111: color_data = 12'b111111111111;
20'b00111011110101011000: color_data = 12'b111111111111;
20'b00111011110101011001: color_data = 12'b111111111111;
20'b00111011110101011010: color_data = 12'b111111111111;
20'b00111011110101011011: color_data = 12'b111111111111;
20'b00111011110101011100: color_data = 12'b111111111111;
20'b00111011110101011101: color_data = 12'b111111111111;
20'b00111011110101011110: color_data = 12'b111111111111;
20'b00111011110101011111: color_data = 12'b111111111111;
20'b00111011110101100000: color_data = 12'b111111111111;
20'b00111011110101100001: color_data = 12'b111111111111;
20'b00111011110101100010: color_data = 12'b111111111111;
20'b00111011110101100011: color_data = 12'b111111111111;
20'b00111011110101100100: color_data = 12'b111111111111;
20'b00111011110101100101: color_data = 12'b111111111111;
20'b00111011110101100110: color_data = 12'b111111111111;
20'b00111011110101100111: color_data = 12'b111111111111;
20'b00111011110101101000: color_data = 12'b111111111111;
20'b00111011110101101001: color_data = 12'b111111111111;
20'b00111011110101101111: color_data = 12'b111111111111;
20'b00111011110101110000: color_data = 12'b111111111111;
20'b00111011110101110001: color_data = 12'b111111111111;
20'b00111011110101110010: color_data = 12'b111111111111;
20'b00111011110101110011: color_data = 12'b111111111111;
20'b00111011110110001101: color_data = 12'b111111111111;
20'b00111011110110001110: color_data = 12'b111111111111;
20'b00111011110110001111: color_data = 12'b111111111111;
20'b00111011110110010000: color_data = 12'b111111111111;
20'b00111011110110010001: color_data = 12'b111111111111;
20'b00111011110110010010: color_data = 12'b111111111111;
20'b00111011110110010011: color_data = 12'b111111111111;
20'b00111011110110010100: color_data = 12'b111111111111;
20'b00111011110110010101: color_data = 12'b111111111111;
20'b00111011110110010110: color_data = 12'b111111111111;
20'b00111011110110010111: color_data = 12'b111111111111;
20'b00111011110110011000: color_data = 12'b111111111111;
20'b00111011110110011001: color_data = 12'b111111111111;
20'b00111011110110011010: color_data = 12'b111111111111;
20'b00111011110110011011: color_data = 12'b111111111111;
20'b00111011110110011100: color_data = 12'b111111111111;
20'b00111011110110011101: color_data = 12'b111111111111;
20'b00111011110110011110: color_data = 12'b111111111111;
20'b00111011110110011111: color_data = 12'b111111111111;
20'b00111011110110100000: color_data = 12'b111111111111;
20'b00111100000100001000: color_data = 12'b111111111111;
20'b00111100000100001001: color_data = 12'b111111111111;
20'b00111100000100001010: color_data = 12'b111111111111;
20'b00111100000100001011: color_data = 12'b111111111111;
20'b00111100000100001100: color_data = 12'b111111111111;
20'b00111100000100100010: color_data = 12'b111111111111;
20'b00111100000100100011: color_data = 12'b111111111111;
20'b00111100000100100100: color_data = 12'b111111111111;
20'b00111100000100100101: color_data = 12'b111111111111;
20'b00111100000100100110: color_data = 12'b111111111111;
20'b00111100000100111100: color_data = 12'b111111111111;
20'b00111100000100111101: color_data = 12'b111111111111;
20'b00111100000100111110: color_data = 12'b111111111111;
20'b00111100000100111111: color_data = 12'b111111111111;
20'b00111100000101000000: color_data = 12'b111111111111;
20'b00111100000101001011: color_data = 12'b111111111111;
20'b00111100000101001100: color_data = 12'b111111111111;
20'b00111100000101001101: color_data = 12'b111111111111;
20'b00111100000101001110: color_data = 12'b111111111111;
20'b00111100000101001111: color_data = 12'b111111111111;
20'b00111100000101010101: color_data = 12'b111111111111;
20'b00111100000101010110: color_data = 12'b111111111111;
20'b00111100000101010111: color_data = 12'b111111111111;
20'b00111100000101011000: color_data = 12'b111111111111;
20'b00111100000101011001: color_data = 12'b111111111111;
20'b00111100000101101111: color_data = 12'b111111111111;
20'b00111100000101110000: color_data = 12'b111111111111;
20'b00111100000101110001: color_data = 12'b111111111111;
20'b00111100000101110010: color_data = 12'b111111111111;
20'b00111100000101110011: color_data = 12'b111111111111;
20'b00111100000110001101: color_data = 12'b111111111111;
20'b00111100000110001110: color_data = 12'b111111111111;
20'b00111100000110001111: color_data = 12'b111111111111;
20'b00111100000110010000: color_data = 12'b111111111111;
20'b00111100000110010001: color_data = 12'b111111111111;
20'b00111100000110010010: color_data = 12'b111111111111;
20'b00111100010100001000: color_data = 12'b111111111111;
20'b00111100010100001001: color_data = 12'b111111111111;
20'b00111100010100001010: color_data = 12'b111111111111;
20'b00111100010100001011: color_data = 12'b111111111111;
20'b00111100010100001100: color_data = 12'b111111111111;
20'b00111100010100100010: color_data = 12'b111111111111;
20'b00111100010100100011: color_data = 12'b111111111111;
20'b00111100010100100100: color_data = 12'b111111111111;
20'b00111100010100100101: color_data = 12'b111111111111;
20'b00111100010100100110: color_data = 12'b111111111111;
20'b00111100010100111100: color_data = 12'b111111111111;
20'b00111100010100111101: color_data = 12'b111111111111;
20'b00111100010100111110: color_data = 12'b111111111111;
20'b00111100010100111111: color_data = 12'b111111111111;
20'b00111100010101000000: color_data = 12'b111111111111;
20'b00111100010101001011: color_data = 12'b111111111111;
20'b00111100010101001100: color_data = 12'b111111111111;
20'b00111100010101001101: color_data = 12'b111111111111;
20'b00111100010101001110: color_data = 12'b111111111111;
20'b00111100010101001111: color_data = 12'b111111111111;
20'b00111100010101010101: color_data = 12'b111111111111;
20'b00111100010101010110: color_data = 12'b111111111111;
20'b00111100010101010111: color_data = 12'b111111111111;
20'b00111100010101011000: color_data = 12'b111111111111;
20'b00111100010101011001: color_data = 12'b111111111111;
20'b00111100010101101111: color_data = 12'b111111111111;
20'b00111100010101110000: color_data = 12'b111111111111;
20'b00111100010101110001: color_data = 12'b111111111111;
20'b00111100010101110010: color_data = 12'b111111111111;
20'b00111100010101110011: color_data = 12'b111111111111;
20'b00111100010110001101: color_data = 12'b111111111111;
20'b00111100010110001110: color_data = 12'b111111111111;
20'b00111100010110001111: color_data = 12'b111111111111;
20'b00111100010110010000: color_data = 12'b111111111111;
20'b00111100010110010001: color_data = 12'b111111111111;
20'b00111100010110010010: color_data = 12'b111111111111;
20'b00111100100100001000: color_data = 12'b111111111111;
20'b00111100100100001001: color_data = 12'b111111111111;
20'b00111100100100001010: color_data = 12'b111111111111;
20'b00111100100100001011: color_data = 12'b111111111111;
20'b00111100100100001100: color_data = 12'b111111111111;
20'b00111100100100100010: color_data = 12'b111111111111;
20'b00111100100100100011: color_data = 12'b111111111111;
20'b00111100100100100100: color_data = 12'b111111111111;
20'b00111100100100100101: color_data = 12'b111111111111;
20'b00111100100100100110: color_data = 12'b111111111111;
20'b00111100100100111100: color_data = 12'b111111111111;
20'b00111100100100111101: color_data = 12'b111111111111;
20'b00111100100100111110: color_data = 12'b111111111111;
20'b00111100100100111111: color_data = 12'b111111111111;
20'b00111100100101000000: color_data = 12'b111111111111;
20'b00111100100101001011: color_data = 12'b111111111111;
20'b00111100100101001100: color_data = 12'b111111111111;
20'b00111100100101001101: color_data = 12'b111111111111;
20'b00111100100101001110: color_data = 12'b111111111111;
20'b00111100100101001111: color_data = 12'b111111111111;
20'b00111100100101010101: color_data = 12'b111111111111;
20'b00111100100101010110: color_data = 12'b111111111111;
20'b00111100100101010111: color_data = 12'b111111111111;
20'b00111100100101011000: color_data = 12'b111111111111;
20'b00111100100101011001: color_data = 12'b111111111111;
20'b00111100100101101111: color_data = 12'b111111111111;
20'b00111100100101110000: color_data = 12'b111111111111;
20'b00111100100101110001: color_data = 12'b111111111111;
20'b00111100100101110010: color_data = 12'b111111111111;
20'b00111100100101110011: color_data = 12'b111111111111;
20'b00111100100110001101: color_data = 12'b111111111111;
20'b00111100100110001110: color_data = 12'b111111111111;
20'b00111100100110001111: color_data = 12'b111111111111;
20'b00111100100110010000: color_data = 12'b111111111111;
20'b00111100100110010001: color_data = 12'b111111111111;
20'b00111100100110010010: color_data = 12'b111111111111;
20'b00111100110100001000: color_data = 12'b111111111111;
20'b00111100110100001001: color_data = 12'b111111111111;
20'b00111100110100001010: color_data = 12'b111111111111;
20'b00111100110100001011: color_data = 12'b111111111111;
20'b00111100110100001100: color_data = 12'b111111111111;
20'b00111100110100100010: color_data = 12'b111111111111;
20'b00111100110100100011: color_data = 12'b111111111111;
20'b00111100110100100100: color_data = 12'b111111111111;
20'b00111100110100100101: color_data = 12'b111111111111;
20'b00111100110100100110: color_data = 12'b111111111111;
20'b00111100110100111100: color_data = 12'b111111111111;
20'b00111100110100111101: color_data = 12'b111111111111;
20'b00111100110100111110: color_data = 12'b111111111111;
20'b00111100110100111111: color_data = 12'b111111111111;
20'b00111100110101000000: color_data = 12'b111111111111;
20'b00111100110101001011: color_data = 12'b111111111111;
20'b00111100110101001100: color_data = 12'b111111111111;
20'b00111100110101001101: color_data = 12'b111111111111;
20'b00111100110101001110: color_data = 12'b111111111111;
20'b00111100110101001111: color_data = 12'b111111111111;
20'b00111100110101010101: color_data = 12'b111111111111;
20'b00111100110101010110: color_data = 12'b111111111111;
20'b00111100110101010111: color_data = 12'b111111111111;
20'b00111100110101011000: color_data = 12'b111111111111;
20'b00111100110101011001: color_data = 12'b111111111111;
20'b00111100110101101111: color_data = 12'b111111111111;
20'b00111100110101110000: color_data = 12'b111111111111;
20'b00111100110101110001: color_data = 12'b111111111111;
20'b00111100110101110010: color_data = 12'b111111111111;
20'b00111100110101110011: color_data = 12'b111111111111;
20'b00111100110110001101: color_data = 12'b111111111111;
20'b00111100110110001110: color_data = 12'b111111111111;
20'b00111100110110001111: color_data = 12'b111111111111;
20'b00111100110110010000: color_data = 12'b111111111111;
20'b00111100110110010001: color_data = 12'b111111111111;
20'b00111100110110010010: color_data = 12'b111111111111;
20'b00111101000100001000: color_data = 12'b111111111111;
20'b00111101000100001001: color_data = 12'b111111111111;
20'b00111101000100001010: color_data = 12'b111111111111;
20'b00111101000100001011: color_data = 12'b111111111111;
20'b00111101000100001100: color_data = 12'b111111111111;
20'b00111101000100001101: color_data = 12'b111111111111;
20'b00111101000100001110: color_data = 12'b111111111111;
20'b00111101000100001111: color_data = 12'b111111111111;
20'b00111101000100010000: color_data = 12'b111111111111;
20'b00111101000100010001: color_data = 12'b111111111111;
20'b00111101000100010010: color_data = 12'b111111111111;
20'b00111101000100010011: color_data = 12'b111111111111;
20'b00111101000100010100: color_data = 12'b111111111111;
20'b00111101000100010101: color_data = 12'b111111111111;
20'b00111101000100010110: color_data = 12'b111111111111;
20'b00111101000100010111: color_data = 12'b111111111111;
20'b00111101000100011000: color_data = 12'b111111111111;
20'b00111101000100011001: color_data = 12'b111111111111;
20'b00111101000100011010: color_data = 12'b111111111111;
20'b00111101000100011011: color_data = 12'b111111111111;
20'b00111101000100011100: color_data = 12'b111111111111;
20'b00111101000100100010: color_data = 12'b111111111111;
20'b00111101000100100011: color_data = 12'b111111111111;
20'b00111101000100100100: color_data = 12'b111111111111;
20'b00111101000100100101: color_data = 12'b111111111111;
20'b00111101000100100110: color_data = 12'b111111111111;
20'b00111101000100100111: color_data = 12'b111111111111;
20'b00111101000100101000: color_data = 12'b111111111111;
20'b00111101000100101001: color_data = 12'b111111111111;
20'b00111101000100101010: color_data = 12'b111111111111;
20'b00111101000100101011: color_data = 12'b111111111111;
20'b00111101000100101100: color_data = 12'b111111111111;
20'b00111101000100101101: color_data = 12'b111111111111;
20'b00111101000100101110: color_data = 12'b111111111111;
20'b00111101000100101111: color_data = 12'b111111111111;
20'b00111101000100110000: color_data = 12'b111111111111;
20'b00111101000100110001: color_data = 12'b111111111111;
20'b00111101000100110010: color_data = 12'b111111111111;
20'b00111101000100110011: color_data = 12'b111111111111;
20'b00111101000100110100: color_data = 12'b111111111111;
20'b00111101000100110101: color_data = 12'b111111111111;
20'b00111101000100111100: color_data = 12'b111111111111;
20'b00111101000100111101: color_data = 12'b111111111111;
20'b00111101000100111110: color_data = 12'b111111111111;
20'b00111101000100111111: color_data = 12'b111111111111;
20'b00111101000101000000: color_data = 12'b111111111111;
20'b00111101000101000001: color_data = 12'b111111111111;
20'b00111101000101000010: color_data = 12'b111111111111;
20'b00111101000101000011: color_data = 12'b111111111111;
20'b00111101000101000100: color_data = 12'b111111111111;
20'b00111101000101000101: color_data = 12'b111111111111;
20'b00111101000101000110: color_data = 12'b111111111111;
20'b00111101000101000111: color_data = 12'b111111111111;
20'b00111101000101001000: color_data = 12'b111111111111;
20'b00111101000101001001: color_data = 12'b111111111111;
20'b00111101000101001010: color_data = 12'b111111111111;
20'b00111101000101010101: color_data = 12'b111111111111;
20'b00111101000101010110: color_data = 12'b111111111111;
20'b00111101000101010111: color_data = 12'b111111111111;
20'b00111101000101011000: color_data = 12'b111111111111;
20'b00111101000101011001: color_data = 12'b111111111111;
20'b00111101000101011010: color_data = 12'b111111111111;
20'b00111101000101011011: color_data = 12'b111111111111;
20'b00111101000101011100: color_data = 12'b111111111111;
20'b00111101000101011101: color_data = 12'b111111111111;
20'b00111101000101011110: color_data = 12'b111111111111;
20'b00111101000101011111: color_data = 12'b111111111111;
20'b00111101000101100000: color_data = 12'b111111111111;
20'b00111101000101100001: color_data = 12'b111111111111;
20'b00111101000101100010: color_data = 12'b111111111111;
20'b00111101000101100011: color_data = 12'b111111111111;
20'b00111101000101100100: color_data = 12'b111111111111;
20'b00111101000101100101: color_data = 12'b111111111111;
20'b00111101000101100110: color_data = 12'b111111111111;
20'b00111101000101100111: color_data = 12'b111111111111;
20'b00111101000101101000: color_data = 12'b111111111111;
20'b00111101000101101001: color_data = 12'b111111111111;
20'b00111101000101101111: color_data = 12'b111111111111;
20'b00111101000101110000: color_data = 12'b111111111111;
20'b00111101000101110001: color_data = 12'b111111111111;
20'b00111101000101110010: color_data = 12'b111111111111;
20'b00111101000101110011: color_data = 12'b111111111111;
20'b00111101000101110100: color_data = 12'b111111111111;
20'b00111101000101110101: color_data = 12'b111111111111;
20'b00111101000101110110: color_data = 12'b111111111111;
20'b00111101000101110111: color_data = 12'b111111111111;
20'b00111101000101111000: color_data = 12'b111111111111;
20'b00111101000101111001: color_data = 12'b111111111111;
20'b00111101000101111010: color_data = 12'b111111111111;
20'b00111101000101111011: color_data = 12'b111111111111;
20'b00111101000101111100: color_data = 12'b111111111111;
20'b00111101000101111101: color_data = 12'b111111111111;
20'b00111101000101111110: color_data = 12'b111111111111;
20'b00111101000101111111: color_data = 12'b111111111111;
20'b00111101000110000000: color_data = 12'b111111111111;
20'b00111101000110000001: color_data = 12'b111111111111;
20'b00111101000110000010: color_data = 12'b111111111111;
20'b00111101000110001101: color_data = 12'b111111111111;
20'b00111101000110001110: color_data = 12'b111111111111;
20'b00111101000110001111: color_data = 12'b111111111111;
20'b00111101000110010000: color_data = 12'b111111111111;
20'b00111101000110010001: color_data = 12'b111111111111;
20'b00111101000110010010: color_data = 12'b111111111111;
20'b00111101000110010011: color_data = 12'b111111111111;
20'b00111101000110010100: color_data = 12'b111111111111;
20'b00111101000110010101: color_data = 12'b111111111111;
20'b00111101000110010110: color_data = 12'b111111111111;
20'b00111101000110010111: color_data = 12'b111111111111;
20'b00111101000110011000: color_data = 12'b111111111111;
20'b00111101000110011001: color_data = 12'b111111111111;
20'b00111101000110011010: color_data = 12'b111111111111;
20'b00111101000110011011: color_data = 12'b111111111111;
20'b00111101000110011100: color_data = 12'b111111111111;
20'b00111101000110011101: color_data = 12'b111111111111;
20'b00111101000110011110: color_data = 12'b111111111111;
20'b00111101000110011111: color_data = 12'b111111111111;
20'b00111101000110100000: color_data = 12'b111111111111;
20'b00111101010100001000: color_data = 12'b111111111111;
20'b00111101010100001001: color_data = 12'b111111111111;
20'b00111101010100001010: color_data = 12'b111111111111;
20'b00111101010100001011: color_data = 12'b111111111111;
20'b00111101010100001100: color_data = 12'b111111111111;
20'b00111101010100001101: color_data = 12'b111111111111;
20'b00111101010100001110: color_data = 12'b111111111111;
20'b00111101010100001111: color_data = 12'b111111111111;
20'b00111101010100010000: color_data = 12'b111111111111;
20'b00111101010100010001: color_data = 12'b111111111111;
20'b00111101010100010010: color_data = 12'b111111111111;
20'b00111101010100010011: color_data = 12'b111111111111;
20'b00111101010100010100: color_data = 12'b111111111111;
20'b00111101010100010101: color_data = 12'b111111111111;
20'b00111101010100010110: color_data = 12'b111111111111;
20'b00111101010100010111: color_data = 12'b111111111111;
20'b00111101010100011000: color_data = 12'b111111111111;
20'b00111101010100011001: color_data = 12'b111111111111;
20'b00111101010100011010: color_data = 12'b111111111111;
20'b00111101010100011011: color_data = 12'b111111111111;
20'b00111101010100011100: color_data = 12'b111111111111;
20'b00111101010100100010: color_data = 12'b111111111111;
20'b00111101010100100011: color_data = 12'b111111111111;
20'b00111101010100100100: color_data = 12'b111111111111;
20'b00111101010100100101: color_data = 12'b111111111111;
20'b00111101010100100110: color_data = 12'b111111111111;
20'b00111101010100100111: color_data = 12'b111111111111;
20'b00111101010100101000: color_data = 12'b111111111111;
20'b00111101010100101001: color_data = 12'b111111111111;
20'b00111101010100101010: color_data = 12'b111111111111;
20'b00111101010100101011: color_data = 12'b111111111111;
20'b00111101010100101100: color_data = 12'b111111111111;
20'b00111101010100101101: color_data = 12'b111111111111;
20'b00111101010100101110: color_data = 12'b111111111111;
20'b00111101010100101111: color_data = 12'b111111111111;
20'b00111101010100110000: color_data = 12'b111111111111;
20'b00111101010100110001: color_data = 12'b111111111111;
20'b00111101010100110010: color_data = 12'b111111111111;
20'b00111101010100110011: color_data = 12'b111111111111;
20'b00111101010100110100: color_data = 12'b111111111111;
20'b00111101010100110101: color_data = 12'b111111111111;
20'b00111101010100111100: color_data = 12'b111111111111;
20'b00111101010100111101: color_data = 12'b111111111111;
20'b00111101010100111110: color_data = 12'b111111111111;
20'b00111101010100111111: color_data = 12'b111111111111;
20'b00111101010101000000: color_data = 12'b111111111111;
20'b00111101010101000001: color_data = 12'b111111111111;
20'b00111101010101000010: color_data = 12'b111111111111;
20'b00111101010101000011: color_data = 12'b111111111111;
20'b00111101010101000100: color_data = 12'b111111111111;
20'b00111101010101000101: color_data = 12'b111111111111;
20'b00111101010101000110: color_data = 12'b111111111111;
20'b00111101010101000111: color_data = 12'b111111111111;
20'b00111101010101001000: color_data = 12'b111111111111;
20'b00111101010101001001: color_data = 12'b111111111111;
20'b00111101010101001010: color_data = 12'b111111111111;
20'b00111101010101010101: color_data = 12'b111111111111;
20'b00111101010101010110: color_data = 12'b111111111111;
20'b00111101010101010111: color_data = 12'b111111111111;
20'b00111101010101011000: color_data = 12'b111111111111;
20'b00111101010101011001: color_data = 12'b111111111111;
20'b00111101010101011010: color_data = 12'b111111111111;
20'b00111101010101011011: color_data = 12'b111111111111;
20'b00111101010101011100: color_data = 12'b111111111111;
20'b00111101010101011101: color_data = 12'b111111111111;
20'b00111101010101011110: color_data = 12'b111111111111;
20'b00111101010101011111: color_data = 12'b111111111111;
20'b00111101010101100000: color_data = 12'b111111111111;
20'b00111101010101100001: color_data = 12'b111111111111;
20'b00111101010101100010: color_data = 12'b111111111111;
20'b00111101010101100011: color_data = 12'b111111111111;
20'b00111101010101100100: color_data = 12'b111111111111;
20'b00111101010101100101: color_data = 12'b111111111111;
20'b00111101010101100110: color_data = 12'b111111111111;
20'b00111101010101100111: color_data = 12'b111111111111;
20'b00111101010101101000: color_data = 12'b111111111111;
20'b00111101010101101001: color_data = 12'b111111111111;
20'b00111101010101101111: color_data = 12'b111111111111;
20'b00111101010101110000: color_data = 12'b111111111111;
20'b00111101010101110001: color_data = 12'b111111111111;
20'b00111101010101110010: color_data = 12'b111111111111;
20'b00111101010101110011: color_data = 12'b111111111111;
20'b00111101010101110100: color_data = 12'b111111111111;
20'b00111101010101110101: color_data = 12'b111111111111;
20'b00111101010101110110: color_data = 12'b111111111111;
20'b00111101010101110111: color_data = 12'b111111111111;
20'b00111101010101111000: color_data = 12'b111111111111;
20'b00111101010101111001: color_data = 12'b111111111111;
20'b00111101010101111010: color_data = 12'b111111111111;
20'b00111101010101111011: color_data = 12'b111111111111;
20'b00111101010101111100: color_data = 12'b111111111111;
20'b00111101010101111101: color_data = 12'b111111111111;
20'b00111101010101111110: color_data = 12'b111111111111;
20'b00111101010101111111: color_data = 12'b111111111111;
20'b00111101010110000000: color_data = 12'b111111111111;
20'b00111101010110000001: color_data = 12'b111111111111;
20'b00111101010110000010: color_data = 12'b111111111111;
20'b00111101010110001101: color_data = 12'b111111111111;
20'b00111101010110001110: color_data = 12'b111111111111;
20'b00111101010110001111: color_data = 12'b111111111111;
20'b00111101010110010000: color_data = 12'b111111111111;
20'b00111101010110010001: color_data = 12'b111111111111;
20'b00111101010110010010: color_data = 12'b111111111111;
20'b00111101010110010011: color_data = 12'b111111111111;
20'b00111101010110010100: color_data = 12'b111111111111;
20'b00111101010110010101: color_data = 12'b111111111111;
20'b00111101010110010110: color_data = 12'b111111111111;
20'b00111101010110010111: color_data = 12'b111111111111;
20'b00111101010110011000: color_data = 12'b111111111111;
20'b00111101010110011001: color_data = 12'b111111111111;
20'b00111101010110011010: color_data = 12'b111111111111;
20'b00111101010110011011: color_data = 12'b111111111111;
20'b00111101010110011100: color_data = 12'b111111111111;
20'b00111101010110011101: color_data = 12'b111111111111;
20'b00111101010110011110: color_data = 12'b111111111111;
20'b00111101010110011111: color_data = 12'b111111111111;
20'b00111101010110100000: color_data = 12'b111111111111;
20'b00111101100100001000: color_data = 12'b111111111111;
20'b00111101100100001001: color_data = 12'b111111111111;
20'b00111101100100001010: color_data = 12'b111111111111;
20'b00111101100100001011: color_data = 12'b111111111111;
20'b00111101100100001100: color_data = 12'b111111111111;
20'b00111101100100001101: color_data = 12'b111111111111;
20'b00111101100100001110: color_data = 12'b111111111111;
20'b00111101100100001111: color_data = 12'b111111111111;
20'b00111101100100010000: color_data = 12'b111111111111;
20'b00111101100100010001: color_data = 12'b111111111111;
20'b00111101100100010010: color_data = 12'b111111111111;
20'b00111101100100010011: color_data = 12'b111111111111;
20'b00111101100100010100: color_data = 12'b111111111111;
20'b00111101100100010101: color_data = 12'b111111111111;
20'b00111101100100010110: color_data = 12'b111111111111;
20'b00111101100100010111: color_data = 12'b111111111111;
20'b00111101100100011000: color_data = 12'b111111111111;
20'b00111101100100011001: color_data = 12'b111111111111;
20'b00111101100100011010: color_data = 12'b111111111111;
20'b00111101100100011011: color_data = 12'b111111111111;
20'b00111101100100011100: color_data = 12'b111111111111;
20'b00111101100100100010: color_data = 12'b111111111111;
20'b00111101100100100011: color_data = 12'b111111111111;
20'b00111101100100100100: color_data = 12'b111111111111;
20'b00111101100100100101: color_data = 12'b111111111111;
20'b00111101100100100110: color_data = 12'b111111111111;
20'b00111101100100100111: color_data = 12'b111111111111;
20'b00111101100100101000: color_data = 12'b111111111111;
20'b00111101100100101001: color_data = 12'b111111111111;
20'b00111101100100101010: color_data = 12'b111111111111;
20'b00111101100100101011: color_data = 12'b111111111111;
20'b00111101100100101100: color_data = 12'b111111111111;
20'b00111101100100101101: color_data = 12'b111111111111;
20'b00111101100100101110: color_data = 12'b111111111111;
20'b00111101100100101111: color_data = 12'b111111111111;
20'b00111101100100110000: color_data = 12'b111111111111;
20'b00111101100100110001: color_data = 12'b111111111111;
20'b00111101100100110010: color_data = 12'b111111111111;
20'b00111101100100110011: color_data = 12'b111111111111;
20'b00111101100100110100: color_data = 12'b111111111111;
20'b00111101100100110101: color_data = 12'b111111111111;
20'b00111101100100111100: color_data = 12'b111111111111;
20'b00111101100100111101: color_data = 12'b111111111111;
20'b00111101100100111110: color_data = 12'b111111111111;
20'b00111101100100111111: color_data = 12'b111111111111;
20'b00111101100101000000: color_data = 12'b111111111111;
20'b00111101100101000001: color_data = 12'b111111111111;
20'b00111101100101000010: color_data = 12'b111111111111;
20'b00111101100101000011: color_data = 12'b111111111111;
20'b00111101100101000100: color_data = 12'b111111111111;
20'b00111101100101000101: color_data = 12'b111111111111;
20'b00111101100101000110: color_data = 12'b111111111111;
20'b00111101100101000111: color_data = 12'b111111111111;
20'b00111101100101001000: color_data = 12'b111111111111;
20'b00111101100101001001: color_data = 12'b111111111111;
20'b00111101100101001010: color_data = 12'b111111111111;
20'b00111101100101010101: color_data = 12'b111111111111;
20'b00111101100101010110: color_data = 12'b111111111111;
20'b00111101100101010111: color_data = 12'b111111111111;
20'b00111101100101011000: color_data = 12'b111111111111;
20'b00111101100101011001: color_data = 12'b111111111111;
20'b00111101100101011010: color_data = 12'b111111111111;
20'b00111101100101011011: color_data = 12'b111111111111;
20'b00111101100101011100: color_data = 12'b111111111111;
20'b00111101100101011101: color_data = 12'b111111111111;
20'b00111101100101011110: color_data = 12'b111111111111;
20'b00111101100101011111: color_data = 12'b111111111111;
20'b00111101100101100000: color_data = 12'b111111111111;
20'b00111101100101100001: color_data = 12'b111111111111;
20'b00111101100101100010: color_data = 12'b111111111111;
20'b00111101100101100011: color_data = 12'b111111111111;
20'b00111101100101100100: color_data = 12'b111111111111;
20'b00111101100101100101: color_data = 12'b111111111111;
20'b00111101100101100110: color_data = 12'b111111111111;
20'b00111101100101100111: color_data = 12'b111111111111;
20'b00111101100101101000: color_data = 12'b111111111111;
20'b00111101100101101001: color_data = 12'b111111111111;
20'b00111101100101101111: color_data = 12'b111111111111;
20'b00111101100101110000: color_data = 12'b111111111111;
20'b00111101100101110001: color_data = 12'b111111111111;
20'b00111101100101110010: color_data = 12'b111111111111;
20'b00111101100101110011: color_data = 12'b111111111111;
20'b00111101100101110100: color_data = 12'b111111111111;
20'b00111101100101110101: color_data = 12'b111111111111;
20'b00111101100101110110: color_data = 12'b111111111111;
20'b00111101100101110111: color_data = 12'b111111111111;
20'b00111101100101111000: color_data = 12'b111111111111;
20'b00111101100101111001: color_data = 12'b111111111111;
20'b00111101100101111010: color_data = 12'b111111111111;
20'b00111101100101111011: color_data = 12'b111111111111;
20'b00111101100101111100: color_data = 12'b111111111111;
20'b00111101100101111101: color_data = 12'b111111111111;
20'b00111101100101111110: color_data = 12'b111111111111;
20'b00111101100101111111: color_data = 12'b111111111111;
20'b00111101100110000000: color_data = 12'b111111111111;
20'b00111101100110000001: color_data = 12'b111111111111;
20'b00111101100110000010: color_data = 12'b111111111111;
20'b00111101100110001101: color_data = 12'b111111111111;
20'b00111101100110001110: color_data = 12'b111111111111;
20'b00111101100110001111: color_data = 12'b111111111111;
20'b00111101100110010000: color_data = 12'b111111111111;
20'b00111101100110010001: color_data = 12'b111111111111;
20'b00111101100110010010: color_data = 12'b111111111111;
20'b00111101100110010011: color_data = 12'b111111111111;
20'b00111101100110010100: color_data = 12'b111111111111;
20'b00111101100110010101: color_data = 12'b111111111111;
20'b00111101100110010110: color_data = 12'b111111111111;
20'b00111101100110010111: color_data = 12'b111111111111;
20'b00111101100110011000: color_data = 12'b111111111111;
20'b00111101100110011001: color_data = 12'b111111111111;
20'b00111101100110011010: color_data = 12'b111111111111;
20'b00111101100110011011: color_data = 12'b111111111111;
20'b00111101100110011100: color_data = 12'b111111111111;
20'b00111101100110011101: color_data = 12'b111111111111;
20'b00111101100110011110: color_data = 12'b111111111111;
20'b00111101100110011111: color_data = 12'b111111111111;
20'b00111101100110100000: color_data = 12'b111111111111;
20'b00111101110100001000: color_data = 12'b111111111111;
20'b00111101110100001001: color_data = 12'b111111111111;
20'b00111101110100001010: color_data = 12'b111111111111;
20'b00111101110100001011: color_data = 12'b111111111111;
20'b00111101110100001100: color_data = 12'b111111111111;
20'b00111101110100001101: color_data = 12'b111111111111;
20'b00111101110100001110: color_data = 12'b111111111111;
20'b00111101110100001111: color_data = 12'b111111111111;
20'b00111101110100010000: color_data = 12'b111111111111;
20'b00111101110100010001: color_data = 12'b111111111111;
20'b00111101110100010010: color_data = 12'b111111111111;
20'b00111101110100010011: color_data = 12'b111111111111;
20'b00111101110100010100: color_data = 12'b111111111111;
20'b00111101110100010101: color_data = 12'b111111111111;
20'b00111101110100010110: color_data = 12'b111111111111;
20'b00111101110100010111: color_data = 12'b111111111111;
20'b00111101110100011000: color_data = 12'b111111111111;
20'b00111101110100011001: color_data = 12'b111111111111;
20'b00111101110100011010: color_data = 12'b111111111111;
20'b00111101110100011011: color_data = 12'b111111111111;
20'b00111101110100011100: color_data = 12'b111111111111;
20'b00111101110100100010: color_data = 12'b111111111111;
20'b00111101110100100011: color_data = 12'b111111111111;
20'b00111101110100100100: color_data = 12'b111111111111;
20'b00111101110100100101: color_data = 12'b111111111111;
20'b00111101110100100110: color_data = 12'b111111111111;
20'b00111101110100100111: color_data = 12'b111111111111;
20'b00111101110100101000: color_data = 12'b111111111111;
20'b00111101110100101001: color_data = 12'b111111111111;
20'b00111101110100101010: color_data = 12'b111111111111;
20'b00111101110100101011: color_data = 12'b111111111111;
20'b00111101110100101100: color_data = 12'b111111111111;
20'b00111101110100101101: color_data = 12'b111111111111;
20'b00111101110100101110: color_data = 12'b111111111111;
20'b00111101110100101111: color_data = 12'b111111111111;
20'b00111101110100110000: color_data = 12'b111111111111;
20'b00111101110100110001: color_data = 12'b111111111111;
20'b00111101110100110010: color_data = 12'b111111111111;
20'b00111101110100110011: color_data = 12'b111111111111;
20'b00111101110100110100: color_data = 12'b111111111111;
20'b00111101110100110101: color_data = 12'b111111111111;
20'b00111101110100111100: color_data = 12'b111111111111;
20'b00111101110100111101: color_data = 12'b111111111111;
20'b00111101110100111110: color_data = 12'b111111111111;
20'b00111101110100111111: color_data = 12'b111111111111;
20'b00111101110101000000: color_data = 12'b111111111111;
20'b00111101110101000001: color_data = 12'b111111111111;
20'b00111101110101000010: color_data = 12'b111111111111;
20'b00111101110101000011: color_data = 12'b111111111111;
20'b00111101110101000100: color_data = 12'b111111111111;
20'b00111101110101000101: color_data = 12'b111111111111;
20'b00111101110101000110: color_data = 12'b111111111111;
20'b00111101110101000111: color_data = 12'b111111111111;
20'b00111101110101001000: color_data = 12'b111111111111;
20'b00111101110101001001: color_data = 12'b111111111111;
20'b00111101110101001010: color_data = 12'b111111111111;
20'b00111101110101010101: color_data = 12'b111111111111;
20'b00111101110101010110: color_data = 12'b111111111111;
20'b00111101110101010111: color_data = 12'b111111111111;
20'b00111101110101011000: color_data = 12'b111111111111;
20'b00111101110101011001: color_data = 12'b111111111111;
20'b00111101110101011010: color_data = 12'b111111111111;
20'b00111101110101011011: color_data = 12'b111111111111;
20'b00111101110101011100: color_data = 12'b111111111111;
20'b00111101110101011101: color_data = 12'b111111111111;
20'b00111101110101011110: color_data = 12'b111111111111;
20'b00111101110101011111: color_data = 12'b111111111111;
20'b00111101110101100000: color_data = 12'b111111111111;
20'b00111101110101100001: color_data = 12'b111111111111;
20'b00111101110101100010: color_data = 12'b111111111111;
20'b00111101110101100011: color_data = 12'b111111111111;
20'b00111101110101100100: color_data = 12'b111111111111;
20'b00111101110101100101: color_data = 12'b111111111111;
20'b00111101110101100110: color_data = 12'b111111111111;
20'b00111101110101100111: color_data = 12'b111111111111;
20'b00111101110101101000: color_data = 12'b111111111111;
20'b00111101110101101001: color_data = 12'b111111111111;
20'b00111101110101101111: color_data = 12'b111111111111;
20'b00111101110101110000: color_data = 12'b111111111111;
20'b00111101110101110001: color_data = 12'b111111111111;
20'b00111101110101110010: color_data = 12'b111111111111;
20'b00111101110101110011: color_data = 12'b111111111111;
20'b00111101110101110100: color_data = 12'b111111111111;
20'b00111101110101110101: color_data = 12'b111111111111;
20'b00111101110101110110: color_data = 12'b111111111111;
20'b00111101110101110111: color_data = 12'b111111111111;
20'b00111101110101111000: color_data = 12'b111111111111;
20'b00111101110101111001: color_data = 12'b111111111111;
20'b00111101110101111010: color_data = 12'b111111111111;
20'b00111101110101111011: color_data = 12'b111111111111;
20'b00111101110101111100: color_data = 12'b111111111111;
20'b00111101110101111101: color_data = 12'b111111111111;
20'b00111101110101111110: color_data = 12'b111111111111;
20'b00111101110101111111: color_data = 12'b111111111111;
20'b00111101110110000000: color_data = 12'b111111111111;
20'b00111101110110000001: color_data = 12'b111111111111;
20'b00111101110110000010: color_data = 12'b111111111111;
20'b00111101110110001101: color_data = 12'b111111111111;
20'b00111101110110001110: color_data = 12'b111111111111;
20'b00111101110110001111: color_data = 12'b111111111111;
20'b00111101110110010000: color_data = 12'b111111111111;
20'b00111101110110010001: color_data = 12'b111111111111;
20'b00111101110110010010: color_data = 12'b111111111111;
20'b00111101110110010011: color_data = 12'b111111111111;
20'b00111101110110010100: color_data = 12'b111111111111;
20'b00111101110110010101: color_data = 12'b111111111111;
20'b00111101110110010110: color_data = 12'b111111111111;
20'b00111101110110010111: color_data = 12'b111111111111;
20'b00111101110110011000: color_data = 12'b111111111111;
20'b00111101110110011001: color_data = 12'b111111111111;
20'b00111101110110011010: color_data = 12'b111111111111;
20'b00111101110110011011: color_data = 12'b111111111111;
20'b00111101110110011100: color_data = 12'b111111111111;
20'b00111101110110011101: color_data = 12'b111111111111;
20'b00111101110110011110: color_data = 12'b111111111111;
20'b00111101110110011111: color_data = 12'b111111111111;
20'b00111101110110100000: color_data = 12'b111111111111;
20'b01000001100011110011: color_data = 12'b111111111111;
20'b01000001100011110100: color_data = 12'b111111111111;
20'b01000001100011110101: color_data = 12'b111111111111;
20'b01000001100011110110: color_data = 12'b111111111111;
20'b01000001100011110111: color_data = 12'b111111111111;
20'b01000001100011111000: color_data = 12'b111111111111;
20'b01000001100011111001: color_data = 12'b111111111111;
20'b01000001100011111010: color_data = 12'b111111111111;
20'b01000001100100010101: color_data = 12'b111111111111;
20'b01000001100100010110: color_data = 12'b111111111111;
20'b01000001100100010111: color_data = 12'b111111111111;
20'b01000001100100011000: color_data = 12'b111111111111;
20'b01000001100100011001: color_data = 12'b111111111111;
20'b01000001100100011010: color_data = 12'b111111111111;
20'b01000001100100011011: color_data = 12'b111111111111;
20'b01000001100100011100: color_data = 12'b111111111111;
20'b01000001100100011101: color_data = 12'b111111111111;
20'b01000001100100011110: color_data = 12'b111111111111;
20'b01000001100100011111: color_data = 12'b111111111111;
20'b01000001100100100000: color_data = 12'b111111111111;
20'b01000001100100100001: color_data = 12'b111111111111;
20'b01000001100100100010: color_data = 12'b111111111111;
20'b01000001100100100011: color_data = 12'b111111111111;
20'b01000001100100100100: color_data = 12'b111111111111;
20'b01000001100100100101: color_data = 12'b111111111111;
20'b01000001100100100110: color_data = 12'b111111111111;
20'b01000001100100100111: color_data = 12'b111111111111;
20'b01000001100100101000: color_data = 12'b111111111111;
20'b01000001100100101001: color_data = 12'b111111111111;
20'b01000001100100101010: color_data = 12'b111111111111;
20'b01000001100100101011: color_data = 12'b111111111111;
20'b01000001100100101100: color_data = 12'b111111111111;
20'b01000001100100101101: color_data = 12'b111111111111;
20'b01000001100100110100: color_data = 12'b111111111111;
20'b01000001100100110101: color_data = 12'b111111111111;
20'b01000001100100110110: color_data = 12'b111111111111;
20'b01000001100100110111: color_data = 12'b111111111111;
20'b01000001100100111000: color_data = 12'b111111111111;
20'b01000001100100111001: color_data = 12'b111111111111;
20'b01000001100100111010: color_data = 12'b111111111111;
20'b01000001100101001000: color_data = 12'b111111111111;
20'b01000001100101001001: color_data = 12'b111111111111;
20'b01000001100101001010: color_data = 12'b111111111111;
20'b01000001100101001011: color_data = 12'b111111111111;
20'b01000001100101001100: color_data = 12'b111111111111;
20'b01000001100101001101: color_data = 12'b111111111111;
20'b01000001100101010100: color_data = 12'b111111111111;
20'b01000001100101010101: color_data = 12'b111111111111;
20'b01000001100101010110: color_data = 12'b111111111111;
20'b01000001100101010111: color_data = 12'b111111111111;
20'b01000001100101011000: color_data = 12'b111111111111;
20'b01000001100101011001: color_data = 12'b111111111111;
20'b01000001100101011010: color_data = 12'b111111111111;
20'b01000001100101011011: color_data = 12'b111111111111;
20'b01000001100101011100: color_data = 12'b111111111111;
20'b01000001100101011101: color_data = 12'b111111111111;
20'b01000001100101011110: color_data = 12'b111111111111;
20'b01000001100101011111: color_data = 12'b111111111111;
20'b01000001100101100000: color_data = 12'b111111111111;
20'b01000001100101100001: color_data = 12'b111111111111;
20'b01000001100101100010: color_data = 12'b111111111111;
20'b01000001100101100011: color_data = 12'b111111111111;
20'b01000001100101100100: color_data = 12'b111111111111;
20'b01000001100101100101: color_data = 12'b111111111111;
20'b01000001100101100110: color_data = 12'b111111111111;
20'b01000001100101100111: color_data = 12'b111111111111;
20'b01000001100101101000: color_data = 12'b111111111111;
20'b01000001100101101001: color_data = 12'b111111111111;
20'b01000001100101101010: color_data = 12'b111111111111;
20'b01000001100101101011: color_data = 12'b111111111111;
20'b01000001100101101100: color_data = 12'b111111111111;
20'b01000001100101101101: color_data = 12'b111111111111;
20'b01000001100101110100: color_data = 12'b111111111111;
20'b01000001100101110101: color_data = 12'b111111111111;
20'b01000001100101110110: color_data = 12'b111111111111;
20'b01000001100101110111: color_data = 12'b111111111111;
20'b01000001100101111000: color_data = 12'b111111111111;
20'b01000001100101111001: color_data = 12'b111111111111;
20'b01000001100110011010: color_data = 12'b111111111111;
20'b01000001100110011011: color_data = 12'b111111111111;
20'b01000001100110011100: color_data = 12'b111111111111;
20'b01000001100110011101: color_data = 12'b111111111111;
20'b01000001100110011110: color_data = 12'b111111111111;
20'b01000001100110011111: color_data = 12'b111111111111;
20'b01000001100110100000: color_data = 12'b111111111111;
20'b01000001100110100001: color_data = 12'b111111111111;
20'b01000001100110100010: color_data = 12'b111111111111;
20'b01000001100110100011: color_data = 12'b111111111111;
20'b01000001100110100100: color_data = 12'b111111111111;
20'b01000001100110100101: color_data = 12'b111111111111;
20'b01000001100110100110: color_data = 12'b111111111111;
20'b01000001100110100111: color_data = 12'b111111111111;
20'b01000001100110101000: color_data = 12'b111111111111;
20'b01000001100110101001: color_data = 12'b111111111111;
20'b01000001100110101010: color_data = 12'b111111111111;
20'b01000001100110101011: color_data = 12'b111111111111;
20'b01000001100110101100: color_data = 12'b111111111111;
20'b01000001100110101101: color_data = 12'b111111111111;
20'b01000001100110101110: color_data = 12'b111111111111;
20'b01000001100110101111: color_data = 12'b111111111111;
20'b01000001100110110000: color_data = 12'b111111111111;
20'b01000001100110110001: color_data = 12'b111111111111;
20'b01000001100110110010: color_data = 12'b111111111111;
20'b01000001100110110011: color_data = 12'b111111111111;
20'b01000001110011110011: color_data = 12'b111111111111;
20'b01000001110011110100: color_data = 12'b111111111111;
20'b01000001110011110101: color_data = 12'b111111111111;
20'b01000001110011110110: color_data = 12'b111111111111;
20'b01000001110011110111: color_data = 12'b111111111111;
20'b01000001110011111000: color_data = 12'b111111111111;
20'b01000001110011111001: color_data = 12'b111111111111;
20'b01000001110011111010: color_data = 12'b111111111111;
20'b01000001110100010101: color_data = 12'b111111111111;
20'b01000001110100010110: color_data = 12'b111111111111;
20'b01000001110100010111: color_data = 12'b111111111111;
20'b01000001110100011000: color_data = 12'b111111111111;
20'b01000001110100011001: color_data = 12'b111111111111;
20'b01000001110100011010: color_data = 12'b111111111111;
20'b01000001110100011011: color_data = 12'b111111111111;
20'b01000001110100011100: color_data = 12'b111111111111;
20'b01000001110100011101: color_data = 12'b111111111111;
20'b01000001110100011110: color_data = 12'b111111111111;
20'b01000001110100011111: color_data = 12'b111111111111;
20'b01000001110100100000: color_data = 12'b111111111111;
20'b01000001110100100001: color_data = 12'b111111111111;
20'b01000001110100100010: color_data = 12'b111111111111;
20'b01000001110100100011: color_data = 12'b111111111111;
20'b01000001110100100100: color_data = 12'b111111111111;
20'b01000001110100100101: color_data = 12'b111111111111;
20'b01000001110100100110: color_data = 12'b111111111111;
20'b01000001110100100111: color_data = 12'b111111111111;
20'b01000001110100101000: color_data = 12'b111111111111;
20'b01000001110100101001: color_data = 12'b111111111111;
20'b01000001110100101010: color_data = 12'b111111111111;
20'b01000001110100101011: color_data = 12'b111111111111;
20'b01000001110100101100: color_data = 12'b111111111111;
20'b01000001110100101101: color_data = 12'b111111111111;
20'b01000001110100110100: color_data = 12'b111111111111;
20'b01000001110100110101: color_data = 12'b111111111111;
20'b01000001110100110110: color_data = 12'b111111111111;
20'b01000001110100110111: color_data = 12'b111111111111;
20'b01000001110100111000: color_data = 12'b111111111111;
20'b01000001110100111001: color_data = 12'b111111111111;
20'b01000001110100111010: color_data = 12'b111111111111;
20'b01000001110101001000: color_data = 12'b111111111111;
20'b01000001110101001001: color_data = 12'b111111111111;
20'b01000001110101001010: color_data = 12'b111111111111;
20'b01000001110101001011: color_data = 12'b111111111111;
20'b01000001110101001100: color_data = 12'b111111111111;
20'b01000001110101001101: color_data = 12'b111111111111;
20'b01000001110101010100: color_data = 12'b111111111111;
20'b01000001110101010101: color_data = 12'b111111111111;
20'b01000001110101010110: color_data = 12'b111111111111;
20'b01000001110101010111: color_data = 12'b111111111111;
20'b01000001110101011000: color_data = 12'b111111111111;
20'b01000001110101011001: color_data = 12'b111111111111;
20'b01000001110101011010: color_data = 12'b111111111111;
20'b01000001110101011011: color_data = 12'b111111111111;
20'b01000001110101011100: color_data = 12'b111111111111;
20'b01000001110101011101: color_data = 12'b111111111111;
20'b01000001110101011110: color_data = 12'b111111111111;
20'b01000001110101011111: color_data = 12'b111111111111;
20'b01000001110101100000: color_data = 12'b111111111111;
20'b01000001110101100001: color_data = 12'b111111111111;
20'b01000001110101100010: color_data = 12'b111111111111;
20'b01000001110101100011: color_data = 12'b111111111111;
20'b01000001110101100100: color_data = 12'b111111111111;
20'b01000001110101100101: color_data = 12'b111111111111;
20'b01000001110101100110: color_data = 12'b111111111111;
20'b01000001110101100111: color_data = 12'b111111111111;
20'b01000001110101101000: color_data = 12'b111111111111;
20'b01000001110101101001: color_data = 12'b111111111111;
20'b01000001110101101010: color_data = 12'b111111111111;
20'b01000001110101101011: color_data = 12'b111111111111;
20'b01000001110101101100: color_data = 12'b111111111111;
20'b01000001110101101101: color_data = 12'b111111111111;
20'b01000001110101110100: color_data = 12'b111111111111;
20'b01000001110101110101: color_data = 12'b111111111111;
20'b01000001110101110110: color_data = 12'b111111111111;
20'b01000001110101110111: color_data = 12'b111111111111;
20'b01000001110101111000: color_data = 12'b111111111111;
20'b01000001110101111001: color_data = 12'b111111111111;
20'b01000001110110011010: color_data = 12'b111111111111;
20'b01000001110110011011: color_data = 12'b111111111111;
20'b01000001110110011100: color_data = 12'b111111111111;
20'b01000001110110011101: color_data = 12'b111111111111;
20'b01000001110110011110: color_data = 12'b111111111111;
20'b01000001110110011111: color_data = 12'b111111111111;
20'b01000001110110100000: color_data = 12'b111111111111;
20'b01000001110110100001: color_data = 12'b111111111111;
20'b01000001110110100010: color_data = 12'b111111111111;
20'b01000001110110100011: color_data = 12'b111111111111;
20'b01000001110110100100: color_data = 12'b111111111111;
20'b01000001110110100101: color_data = 12'b111111111111;
20'b01000001110110100110: color_data = 12'b111111111111;
20'b01000001110110100111: color_data = 12'b111111111111;
20'b01000001110110101000: color_data = 12'b111111111111;
20'b01000001110110101001: color_data = 12'b111111111111;
20'b01000001110110101010: color_data = 12'b111111111111;
20'b01000001110110101011: color_data = 12'b111111111111;
20'b01000001110110101100: color_data = 12'b111111111111;
20'b01000001110110101101: color_data = 12'b111111111111;
20'b01000001110110101110: color_data = 12'b111111111111;
20'b01000001110110101111: color_data = 12'b111111111111;
20'b01000001110110110000: color_data = 12'b111111111111;
20'b01000001110110110001: color_data = 12'b111111111111;
20'b01000001110110110010: color_data = 12'b111111111111;
20'b01000001110110110011: color_data = 12'b111111111111;
20'b01000010000011110011: color_data = 12'b111111111111;
20'b01000010000011110100: color_data = 12'b111111111111;
20'b01000010000011110101: color_data = 12'b111111111111;
20'b01000010000011110110: color_data = 12'b111111111111;
20'b01000010000011110111: color_data = 12'b111111111111;
20'b01000010000011111000: color_data = 12'b111111111111;
20'b01000010000011111001: color_data = 12'b111111111111;
20'b01000010000011111010: color_data = 12'b111111111111;
20'b01000010000100010101: color_data = 12'b111111111111;
20'b01000010000100010110: color_data = 12'b111111111111;
20'b01000010000100010111: color_data = 12'b111111111111;
20'b01000010000100011000: color_data = 12'b111111111111;
20'b01000010000100011001: color_data = 12'b111111111111;
20'b01000010000100011010: color_data = 12'b111111111111;
20'b01000010000100011011: color_data = 12'b111111111111;
20'b01000010000100011100: color_data = 12'b111111111111;
20'b01000010000100011101: color_data = 12'b111111111111;
20'b01000010000100011110: color_data = 12'b111111111111;
20'b01000010000100011111: color_data = 12'b111111111111;
20'b01000010000100100000: color_data = 12'b111111111111;
20'b01000010000100100001: color_data = 12'b111111111111;
20'b01000010000100100010: color_data = 12'b111111111111;
20'b01000010000100100011: color_data = 12'b111111111111;
20'b01000010000100100100: color_data = 12'b111111111111;
20'b01000010000100100101: color_data = 12'b111111111111;
20'b01000010000100100110: color_data = 12'b111111111111;
20'b01000010000100100111: color_data = 12'b111111111111;
20'b01000010000100101000: color_data = 12'b111111111111;
20'b01000010000100101001: color_data = 12'b111111111111;
20'b01000010000100101010: color_data = 12'b111111111111;
20'b01000010000100101011: color_data = 12'b111111111111;
20'b01000010000100101100: color_data = 12'b111111111111;
20'b01000010000100101101: color_data = 12'b111111111111;
20'b01000010000100110100: color_data = 12'b111111111111;
20'b01000010000100110101: color_data = 12'b111111111111;
20'b01000010000100110110: color_data = 12'b111111111111;
20'b01000010000100110111: color_data = 12'b111111111111;
20'b01000010000100111000: color_data = 12'b111111111111;
20'b01000010000100111001: color_data = 12'b111111111111;
20'b01000010000100111010: color_data = 12'b111111111111;
20'b01000010000101001000: color_data = 12'b111111111111;
20'b01000010000101001001: color_data = 12'b111111111111;
20'b01000010000101001010: color_data = 12'b111111111111;
20'b01000010000101001011: color_data = 12'b111111111111;
20'b01000010000101001100: color_data = 12'b111111111111;
20'b01000010000101001101: color_data = 12'b111111111111;
20'b01000010000101010100: color_data = 12'b111111111111;
20'b01000010000101010101: color_data = 12'b111111111111;
20'b01000010000101010110: color_data = 12'b111111111111;
20'b01000010000101010111: color_data = 12'b111111111111;
20'b01000010000101011000: color_data = 12'b111111111111;
20'b01000010000101011001: color_data = 12'b111111111111;
20'b01000010000101011010: color_data = 12'b111111111111;
20'b01000010000101011011: color_data = 12'b111111111111;
20'b01000010000101011100: color_data = 12'b111111111111;
20'b01000010000101011101: color_data = 12'b111111111111;
20'b01000010000101011110: color_data = 12'b111111111111;
20'b01000010000101011111: color_data = 12'b111111111111;
20'b01000010000101100000: color_data = 12'b111111111111;
20'b01000010000101100001: color_data = 12'b111111111111;
20'b01000010000101100010: color_data = 12'b111111111111;
20'b01000010000101100011: color_data = 12'b111111111111;
20'b01000010000101100100: color_data = 12'b111111111111;
20'b01000010000101100101: color_data = 12'b111111111111;
20'b01000010000101100110: color_data = 12'b111111111111;
20'b01000010000101100111: color_data = 12'b111111111111;
20'b01000010000101101000: color_data = 12'b111111111111;
20'b01000010000101101001: color_data = 12'b111111111111;
20'b01000010000101101010: color_data = 12'b111111111111;
20'b01000010000101101011: color_data = 12'b111111111111;
20'b01000010000101101100: color_data = 12'b111111111111;
20'b01000010000101101101: color_data = 12'b111111111111;
20'b01000010000101110100: color_data = 12'b111111111111;
20'b01000010000101110101: color_data = 12'b111111111111;
20'b01000010000101110110: color_data = 12'b111111111111;
20'b01000010000101110111: color_data = 12'b111111111111;
20'b01000010000101111000: color_data = 12'b111111111111;
20'b01000010000101111001: color_data = 12'b111111111111;
20'b01000010000110011010: color_data = 12'b111111111111;
20'b01000010000110011011: color_data = 12'b111111111111;
20'b01000010000110011100: color_data = 12'b111111111111;
20'b01000010000110011101: color_data = 12'b111111111111;
20'b01000010000110011110: color_data = 12'b111111111111;
20'b01000010000110011111: color_data = 12'b111111111111;
20'b01000010000110100000: color_data = 12'b111111111111;
20'b01000010000110100001: color_data = 12'b111111111111;
20'b01000010000110100010: color_data = 12'b111111111111;
20'b01000010000110100011: color_data = 12'b111111111111;
20'b01000010000110100100: color_data = 12'b111111111111;
20'b01000010000110100101: color_data = 12'b111111111111;
20'b01000010000110100110: color_data = 12'b111111111111;
20'b01000010000110100111: color_data = 12'b111111111111;
20'b01000010000110101000: color_data = 12'b111111111111;
20'b01000010000110101001: color_data = 12'b111111111111;
20'b01000010000110101010: color_data = 12'b111111111111;
20'b01000010000110101011: color_data = 12'b111111111111;
20'b01000010000110101100: color_data = 12'b111111111111;
20'b01000010000110101101: color_data = 12'b111111111111;
20'b01000010000110101110: color_data = 12'b111111111111;
20'b01000010000110101111: color_data = 12'b111111111111;
20'b01000010000110110000: color_data = 12'b111111111111;
20'b01000010000110110001: color_data = 12'b111111111111;
20'b01000010000110110010: color_data = 12'b111111111111;
20'b01000010000110110011: color_data = 12'b111111111111;
20'b01000010010011110011: color_data = 12'b111111111111;
20'b01000010010011110100: color_data = 12'b111111111111;
20'b01000010010011110101: color_data = 12'b111111111111;
20'b01000010010011110110: color_data = 12'b111111111111;
20'b01000010010011110111: color_data = 12'b111111111111;
20'b01000010010011111000: color_data = 12'b111111111111;
20'b01000010010011111001: color_data = 12'b111111111111;
20'b01000010010011111010: color_data = 12'b111111111111;
20'b01000010010100010101: color_data = 12'b111111111111;
20'b01000010010100010110: color_data = 12'b111111111111;
20'b01000010010100010111: color_data = 12'b111111111111;
20'b01000010010100011000: color_data = 12'b111111111111;
20'b01000010010100011001: color_data = 12'b111111111111;
20'b01000010010100011010: color_data = 12'b111111111111;
20'b01000010010100011011: color_data = 12'b111111111111;
20'b01000010010100011100: color_data = 12'b111111111111;
20'b01000010010100011101: color_data = 12'b111111111111;
20'b01000010010100011110: color_data = 12'b111111111111;
20'b01000010010100011111: color_data = 12'b111111111111;
20'b01000010010100100000: color_data = 12'b111111111111;
20'b01000010010100100001: color_data = 12'b111111111111;
20'b01000010010100100010: color_data = 12'b111111111111;
20'b01000010010100100011: color_data = 12'b111111111111;
20'b01000010010100100100: color_data = 12'b111111111111;
20'b01000010010100100101: color_data = 12'b111111111111;
20'b01000010010100100110: color_data = 12'b111111111111;
20'b01000010010100100111: color_data = 12'b111111111111;
20'b01000010010100101000: color_data = 12'b111111111111;
20'b01000010010100101001: color_data = 12'b111111111111;
20'b01000010010100101010: color_data = 12'b111111111111;
20'b01000010010100101011: color_data = 12'b111111111111;
20'b01000010010100101100: color_data = 12'b111111111111;
20'b01000010010100101101: color_data = 12'b111111111111;
20'b01000010010100110100: color_data = 12'b111111111111;
20'b01000010010100110101: color_data = 12'b111111111111;
20'b01000010010100110110: color_data = 12'b111111111111;
20'b01000010010100110111: color_data = 12'b111111111111;
20'b01000010010100111000: color_data = 12'b111111111111;
20'b01000010010100111001: color_data = 12'b111111111111;
20'b01000010010100111010: color_data = 12'b111111111111;
20'b01000010010101001000: color_data = 12'b111111111111;
20'b01000010010101001001: color_data = 12'b111111111111;
20'b01000010010101001010: color_data = 12'b111111111111;
20'b01000010010101001011: color_data = 12'b111111111111;
20'b01000010010101001100: color_data = 12'b111111111111;
20'b01000010010101001101: color_data = 12'b111111111111;
20'b01000010010101010100: color_data = 12'b111111111111;
20'b01000010010101010101: color_data = 12'b111111111111;
20'b01000010010101010110: color_data = 12'b111111111111;
20'b01000010010101010111: color_data = 12'b111111111111;
20'b01000010010101011000: color_data = 12'b111111111111;
20'b01000010010101011001: color_data = 12'b111111111111;
20'b01000010010101011010: color_data = 12'b111111111111;
20'b01000010010101011011: color_data = 12'b111111111111;
20'b01000010010101011100: color_data = 12'b111111111111;
20'b01000010010101011101: color_data = 12'b111111111111;
20'b01000010010101011110: color_data = 12'b111111111111;
20'b01000010010101011111: color_data = 12'b111111111111;
20'b01000010010101100000: color_data = 12'b111111111111;
20'b01000010010101100001: color_data = 12'b111111111111;
20'b01000010010101100010: color_data = 12'b111111111111;
20'b01000010010101100011: color_data = 12'b111111111111;
20'b01000010010101100100: color_data = 12'b111111111111;
20'b01000010010101100101: color_data = 12'b111111111111;
20'b01000010010101100110: color_data = 12'b111111111111;
20'b01000010010101100111: color_data = 12'b111111111111;
20'b01000010010101101000: color_data = 12'b111111111111;
20'b01000010010101101001: color_data = 12'b111111111111;
20'b01000010010101101010: color_data = 12'b111111111111;
20'b01000010010101101011: color_data = 12'b111111111111;
20'b01000010010101101100: color_data = 12'b111111111111;
20'b01000010010101101101: color_data = 12'b111111111111;
20'b01000010010101110100: color_data = 12'b111111111111;
20'b01000010010101110101: color_data = 12'b111111111111;
20'b01000010010101110110: color_data = 12'b111111111111;
20'b01000010010101110111: color_data = 12'b111111111111;
20'b01000010010101111000: color_data = 12'b111111111111;
20'b01000010010101111001: color_data = 12'b111111111111;
20'b01000010010110011010: color_data = 12'b111111111111;
20'b01000010010110011011: color_data = 12'b111111111111;
20'b01000010010110011100: color_data = 12'b111111111111;
20'b01000010010110011101: color_data = 12'b111111111111;
20'b01000010010110011110: color_data = 12'b111111111111;
20'b01000010010110011111: color_data = 12'b111111111111;
20'b01000010010110100000: color_data = 12'b111111111111;
20'b01000010010110100001: color_data = 12'b111111111111;
20'b01000010010110100010: color_data = 12'b111111111111;
20'b01000010010110100011: color_data = 12'b111111111111;
20'b01000010010110100100: color_data = 12'b111111111111;
20'b01000010010110100101: color_data = 12'b111111111111;
20'b01000010010110100110: color_data = 12'b111111111111;
20'b01000010010110100111: color_data = 12'b111111111111;
20'b01000010010110101000: color_data = 12'b111111111111;
20'b01000010010110101001: color_data = 12'b111111111111;
20'b01000010010110101010: color_data = 12'b111111111111;
20'b01000010010110101011: color_data = 12'b111111111111;
20'b01000010010110101100: color_data = 12'b111111111111;
20'b01000010010110101101: color_data = 12'b111111111111;
20'b01000010010110101110: color_data = 12'b111111111111;
20'b01000010010110101111: color_data = 12'b111111111111;
20'b01000010010110110000: color_data = 12'b111111111111;
20'b01000010010110110001: color_data = 12'b111111111111;
20'b01000010010110110010: color_data = 12'b111111111111;
20'b01000010010110110011: color_data = 12'b111111111111;
20'b01000010100011110011: color_data = 12'b111111111111;
20'b01000010100011110100: color_data = 12'b111111111111;
20'b01000010100011110101: color_data = 12'b111111111111;
20'b01000010100011110110: color_data = 12'b111111111111;
20'b01000010100011110111: color_data = 12'b111111111111;
20'b01000010100011111000: color_data = 12'b111111111111;
20'b01000010100011111001: color_data = 12'b111111111111;
20'b01000010100011111010: color_data = 12'b111111111111;
20'b01000010100100010101: color_data = 12'b111111111111;
20'b01000010100100010110: color_data = 12'b111111111111;
20'b01000010100100010111: color_data = 12'b111111111111;
20'b01000010100100011000: color_data = 12'b111111111111;
20'b01000010100100011001: color_data = 12'b111111111111;
20'b01000010100100011010: color_data = 12'b111111111111;
20'b01000010100100011011: color_data = 12'b111111111111;
20'b01000010100100011100: color_data = 12'b111111111111;
20'b01000010100100011101: color_data = 12'b111111111111;
20'b01000010100100011110: color_data = 12'b111111111111;
20'b01000010100100011111: color_data = 12'b111111111111;
20'b01000010100100100000: color_data = 12'b111111111111;
20'b01000010100100100001: color_data = 12'b111111111111;
20'b01000010100100100010: color_data = 12'b111111111111;
20'b01000010100100100011: color_data = 12'b111111111111;
20'b01000010100100100100: color_data = 12'b111111111111;
20'b01000010100100100101: color_data = 12'b111111111111;
20'b01000010100100100110: color_data = 12'b111111111111;
20'b01000010100100100111: color_data = 12'b111111111111;
20'b01000010100100101000: color_data = 12'b111111111111;
20'b01000010100100101001: color_data = 12'b111111111111;
20'b01000010100100101010: color_data = 12'b111111111111;
20'b01000010100100101011: color_data = 12'b111111111111;
20'b01000010100100101100: color_data = 12'b111111111111;
20'b01000010100100101101: color_data = 12'b111111111111;
20'b01000010100100110100: color_data = 12'b111111111111;
20'b01000010100100110101: color_data = 12'b111111111111;
20'b01000010100100110110: color_data = 12'b111111111111;
20'b01000010100100110111: color_data = 12'b111111111111;
20'b01000010100100111000: color_data = 12'b111111111111;
20'b01000010100100111001: color_data = 12'b111111111111;
20'b01000010100100111010: color_data = 12'b111111111111;
20'b01000010100101001000: color_data = 12'b111111111111;
20'b01000010100101001001: color_data = 12'b111111111111;
20'b01000010100101001010: color_data = 12'b111111111111;
20'b01000010100101001011: color_data = 12'b111111111111;
20'b01000010100101001100: color_data = 12'b111111111111;
20'b01000010100101001101: color_data = 12'b111111111111;
20'b01000010100101010100: color_data = 12'b111111111111;
20'b01000010100101010101: color_data = 12'b111111111111;
20'b01000010100101010110: color_data = 12'b111111111111;
20'b01000010100101010111: color_data = 12'b111111111111;
20'b01000010100101011000: color_data = 12'b111111111111;
20'b01000010100101011001: color_data = 12'b111111111111;
20'b01000010100101011010: color_data = 12'b111111111111;
20'b01000010100101011011: color_data = 12'b111111111111;
20'b01000010100101011100: color_data = 12'b111111111111;
20'b01000010100101011101: color_data = 12'b111111111111;
20'b01000010100101011110: color_data = 12'b111111111111;
20'b01000010100101011111: color_data = 12'b111111111111;
20'b01000010100101100000: color_data = 12'b111111111111;
20'b01000010100101100001: color_data = 12'b111111111111;
20'b01000010100101100010: color_data = 12'b111111111111;
20'b01000010100101100011: color_data = 12'b111111111111;
20'b01000010100101100100: color_data = 12'b111111111111;
20'b01000010100101100101: color_data = 12'b111111111111;
20'b01000010100101100110: color_data = 12'b111111111111;
20'b01000010100101100111: color_data = 12'b111111111111;
20'b01000010100101101000: color_data = 12'b111111111111;
20'b01000010100101101001: color_data = 12'b111111111111;
20'b01000010100101101010: color_data = 12'b111111111111;
20'b01000010100101101011: color_data = 12'b111111111111;
20'b01000010100101101100: color_data = 12'b111111111111;
20'b01000010100101101101: color_data = 12'b111111111111;
20'b01000010100101110100: color_data = 12'b111111111111;
20'b01000010100101110101: color_data = 12'b111111111111;
20'b01000010100101110110: color_data = 12'b111111111111;
20'b01000010100101110111: color_data = 12'b111111111111;
20'b01000010100101111000: color_data = 12'b111111111111;
20'b01000010100101111001: color_data = 12'b111111111111;
20'b01000010100110011010: color_data = 12'b111111111111;
20'b01000010100110011011: color_data = 12'b111111111111;
20'b01000010100110011100: color_data = 12'b111111111111;
20'b01000010100110011101: color_data = 12'b111111111111;
20'b01000010100110011110: color_data = 12'b111111111111;
20'b01000010100110011111: color_data = 12'b111111111111;
20'b01000010100110100000: color_data = 12'b111111111111;
20'b01000010100110100001: color_data = 12'b111111111111;
20'b01000010100110100010: color_data = 12'b111111111111;
20'b01000010100110100011: color_data = 12'b111111111111;
20'b01000010100110100100: color_data = 12'b111111111111;
20'b01000010100110100101: color_data = 12'b111111111111;
20'b01000010100110100110: color_data = 12'b111111111111;
20'b01000010100110100111: color_data = 12'b111111111111;
20'b01000010100110101000: color_data = 12'b111111111111;
20'b01000010100110101001: color_data = 12'b111111111111;
20'b01000010100110101010: color_data = 12'b111111111111;
20'b01000010100110101011: color_data = 12'b111111111111;
20'b01000010100110101100: color_data = 12'b111111111111;
20'b01000010100110101101: color_data = 12'b111111111111;
20'b01000010100110101110: color_data = 12'b111111111111;
20'b01000010100110101111: color_data = 12'b111111111111;
20'b01000010100110110000: color_data = 12'b111111111111;
20'b01000010100110110001: color_data = 12'b111111111111;
20'b01000010100110110010: color_data = 12'b111111111111;
20'b01000010100110110011: color_data = 12'b111111111111;
20'b01000010110011110011: color_data = 12'b111111111111;
20'b01000010110011110100: color_data = 12'b111111111111;
20'b01000010110011110101: color_data = 12'b111111111111;
20'b01000010110011110110: color_data = 12'b111111111111;
20'b01000010110011110111: color_data = 12'b111111111111;
20'b01000010110011111000: color_data = 12'b111111111111;
20'b01000010110011111001: color_data = 12'b111111111111;
20'b01000010110011111010: color_data = 12'b111111111111;
20'b01000010110100010101: color_data = 12'b111111111111;
20'b01000010110100010110: color_data = 12'b111111111111;
20'b01000010110100010111: color_data = 12'b111111111111;
20'b01000010110100011000: color_data = 12'b111111111111;
20'b01000010110100011001: color_data = 12'b111111111111;
20'b01000010110100011010: color_data = 12'b111111111111;
20'b01000010110100011011: color_data = 12'b111111111111;
20'b01000010110100011100: color_data = 12'b111111111111;
20'b01000010110100011101: color_data = 12'b111111111111;
20'b01000010110100011110: color_data = 12'b111111111111;
20'b01000010110100011111: color_data = 12'b111111111111;
20'b01000010110100100000: color_data = 12'b111111111111;
20'b01000010110100100001: color_data = 12'b111111111111;
20'b01000010110100100010: color_data = 12'b111111111111;
20'b01000010110100100011: color_data = 12'b111111111111;
20'b01000010110100100100: color_data = 12'b111111111111;
20'b01000010110100100101: color_data = 12'b111111111111;
20'b01000010110100100110: color_data = 12'b111111111111;
20'b01000010110100100111: color_data = 12'b111111111111;
20'b01000010110100101000: color_data = 12'b111111111111;
20'b01000010110100101001: color_data = 12'b111111111111;
20'b01000010110100101010: color_data = 12'b111111111111;
20'b01000010110100101011: color_data = 12'b111111111111;
20'b01000010110100101100: color_data = 12'b111111111111;
20'b01000010110100101101: color_data = 12'b111111111111;
20'b01000010110100110100: color_data = 12'b111111111111;
20'b01000010110100110101: color_data = 12'b111111111111;
20'b01000010110100110110: color_data = 12'b111111111111;
20'b01000010110100110111: color_data = 12'b111111111111;
20'b01000010110100111000: color_data = 12'b111111111111;
20'b01000010110100111001: color_data = 12'b111111111111;
20'b01000010110100111010: color_data = 12'b111111111111;
20'b01000010110101001000: color_data = 12'b111111111111;
20'b01000010110101001001: color_data = 12'b111111111111;
20'b01000010110101001010: color_data = 12'b111111111111;
20'b01000010110101001011: color_data = 12'b111111111111;
20'b01000010110101001100: color_data = 12'b111111111111;
20'b01000010110101001101: color_data = 12'b111111111111;
20'b01000010110101010100: color_data = 12'b111111111111;
20'b01000010110101010101: color_data = 12'b111111111111;
20'b01000010110101010110: color_data = 12'b111111111111;
20'b01000010110101010111: color_data = 12'b111111111111;
20'b01000010110101011000: color_data = 12'b111111111111;
20'b01000010110101011001: color_data = 12'b111111111111;
20'b01000010110101011010: color_data = 12'b111111111111;
20'b01000010110101011011: color_data = 12'b111111111111;
20'b01000010110101011100: color_data = 12'b111111111111;
20'b01000010110101011101: color_data = 12'b111111111111;
20'b01000010110101011110: color_data = 12'b111111111111;
20'b01000010110101011111: color_data = 12'b111111111111;
20'b01000010110101100000: color_data = 12'b111111111111;
20'b01000010110101100001: color_data = 12'b111111111111;
20'b01000010110101100010: color_data = 12'b111111111111;
20'b01000010110101100011: color_data = 12'b111111111111;
20'b01000010110101100100: color_data = 12'b111111111111;
20'b01000010110101100101: color_data = 12'b111111111111;
20'b01000010110101100110: color_data = 12'b111111111111;
20'b01000010110101100111: color_data = 12'b111111111111;
20'b01000010110101101000: color_data = 12'b111111111111;
20'b01000010110101101001: color_data = 12'b111111111111;
20'b01000010110101101010: color_data = 12'b111111111111;
20'b01000010110101101011: color_data = 12'b111111111111;
20'b01000010110101101100: color_data = 12'b111111111111;
20'b01000010110101101101: color_data = 12'b111111111111;
20'b01000010110101110100: color_data = 12'b111111111111;
20'b01000010110101110101: color_data = 12'b111111111111;
20'b01000010110101110110: color_data = 12'b111111111111;
20'b01000010110101110111: color_data = 12'b111111111111;
20'b01000010110101111000: color_data = 12'b111111111111;
20'b01000010110101111001: color_data = 12'b111111111111;
20'b01000010110110011010: color_data = 12'b111111111111;
20'b01000010110110011011: color_data = 12'b111111111111;
20'b01000010110110011100: color_data = 12'b111111111111;
20'b01000010110110011101: color_data = 12'b111111111111;
20'b01000010110110011110: color_data = 12'b111111111111;
20'b01000010110110011111: color_data = 12'b111111111111;
20'b01000010110110100000: color_data = 12'b111111111111;
20'b01000010110110100001: color_data = 12'b111111111111;
20'b01000010110110100010: color_data = 12'b111111111111;
20'b01000010110110100011: color_data = 12'b111111111111;
20'b01000010110110100100: color_data = 12'b111111111111;
20'b01000010110110100101: color_data = 12'b111111111111;
20'b01000010110110100110: color_data = 12'b111111111111;
20'b01000010110110100111: color_data = 12'b111111111111;
20'b01000010110110101000: color_data = 12'b111111111111;
20'b01000010110110101001: color_data = 12'b111111111111;
20'b01000010110110101010: color_data = 12'b111111111111;
20'b01000010110110101011: color_data = 12'b111111111111;
20'b01000010110110101100: color_data = 12'b111111111111;
20'b01000010110110101101: color_data = 12'b111111111111;
20'b01000010110110101110: color_data = 12'b111111111111;
20'b01000010110110101111: color_data = 12'b111111111111;
20'b01000010110110110000: color_data = 12'b111111111111;
20'b01000010110110110001: color_data = 12'b111111111111;
20'b01000010110110110010: color_data = 12'b111111111111;
20'b01000010110110110011: color_data = 12'b111111111111;
20'b01000011000011110011: color_data = 12'b111111111111;
20'b01000011000011110100: color_data = 12'b111111111111;
20'b01000011000011110101: color_data = 12'b111111111111;
20'b01000011000011110110: color_data = 12'b111111111111;
20'b01000011000011110111: color_data = 12'b111111111111;
20'b01000011000011111000: color_data = 12'b111111111111;
20'b01000011000011111001: color_data = 12'b111111111111;
20'b01000011000011111010: color_data = 12'b111111111111;
20'b01000011000100010101: color_data = 12'b111111111111;
20'b01000011000100010110: color_data = 12'b111111111111;
20'b01000011000100010111: color_data = 12'b111111111111;
20'b01000011000100011000: color_data = 12'b111111111111;
20'b01000011000100011001: color_data = 12'b111111111111;
20'b01000011000100011010: color_data = 12'b111111111111;
20'b01000011000100110100: color_data = 12'b111111111111;
20'b01000011000100110101: color_data = 12'b111111111111;
20'b01000011000100110110: color_data = 12'b111111111111;
20'b01000011000100110111: color_data = 12'b111111111111;
20'b01000011000100111000: color_data = 12'b111111111111;
20'b01000011000100111001: color_data = 12'b111111111111;
20'b01000011000100111010: color_data = 12'b111111111111;
20'b01000011000101001000: color_data = 12'b111111111111;
20'b01000011000101001001: color_data = 12'b111111111111;
20'b01000011000101001010: color_data = 12'b111111111111;
20'b01000011000101001011: color_data = 12'b111111111111;
20'b01000011000101001100: color_data = 12'b111111111111;
20'b01000011000101001101: color_data = 12'b111111111111;
20'b01000011000101010100: color_data = 12'b111111111111;
20'b01000011000101010101: color_data = 12'b111111111111;
20'b01000011000101010110: color_data = 12'b111111111111;
20'b01000011000101010111: color_data = 12'b111111111111;
20'b01000011000101011000: color_data = 12'b111111111111;
20'b01000011000101011001: color_data = 12'b111111111111;
20'b01000011000101011010: color_data = 12'b111111111111;
20'b01000011000101110100: color_data = 12'b111111111111;
20'b01000011000101110101: color_data = 12'b111111111111;
20'b01000011000101110110: color_data = 12'b111111111111;
20'b01000011000101110111: color_data = 12'b111111111111;
20'b01000011000101111000: color_data = 12'b111111111111;
20'b01000011000101111001: color_data = 12'b111111111111;
20'b01000011000110101101: color_data = 12'b111111111111;
20'b01000011000110101110: color_data = 12'b111111111111;
20'b01000011000110101111: color_data = 12'b111111111111;
20'b01000011000110110000: color_data = 12'b111111111111;
20'b01000011000110110001: color_data = 12'b111111111111;
20'b01000011000110110010: color_data = 12'b111111111111;
20'b01000011000110110011: color_data = 12'b111111111111;
20'b01000011010011110011: color_data = 12'b111111111111;
20'b01000011010011110100: color_data = 12'b111111111111;
20'b01000011010011110101: color_data = 12'b111111111111;
20'b01000011010011110110: color_data = 12'b111111111111;
20'b01000011010011110111: color_data = 12'b111111111111;
20'b01000011010011111000: color_data = 12'b111111111111;
20'b01000011010011111001: color_data = 12'b111111111111;
20'b01000011010011111010: color_data = 12'b111111111111;
20'b01000011010100010101: color_data = 12'b111111111111;
20'b01000011010100010110: color_data = 12'b111111111111;
20'b01000011010100010111: color_data = 12'b111111111111;
20'b01000011010100011000: color_data = 12'b111111111111;
20'b01000011010100011001: color_data = 12'b111111111111;
20'b01000011010100011010: color_data = 12'b111111111111;
20'b01000011010100110100: color_data = 12'b111111111111;
20'b01000011010100110101: color_data = 12'b111111111111;
20'b01000011010100110110: color_data = 12'b111111111111;
20'b01000011010100110111: color_data = 12'b111111111111;
20'b01000011010100111000: color_data = 12'b111111111111;
20'b01000011010100111001: color_data = 12'b111111111111;
20'b01000011010100111010: color_data = 12'b111111111111;
20'b01000011010101001000: color_data = 12'b111111111111;
20'b01000011010101001001: color_data = 12'b111111111111;
20'b01000011010101001010: color_data = 12'b111111111111;
20'b01000011010101001011: color_data = 12'b111111111111;
20'b01000011010101001100: color_data = 12'b111111111111;
20'b01000011010101001101: color_data = 12'b111111111111;
20'b01000011010101010100: color_data = 12'b111111111111;
20'b01000011010101010101: color_data = 12'b111111111111;
20'b01000011010101010110: color_data = 12'b111111111111;
20'b01000011010101010111: color_data = 12'b111111111111;
20'b01000011010101011000: color_data = 12'b111111111111;
20'b01000011010101011001: color_data = 12'b111111111111;
20'b01000011010101011010: color_data = 12'b111111111111;
20'b01000011010101110100: color_data = 12'b111111111111;
20'b01000011010101110101: color_data = 12'b111111111111;
20'b01000011010101110110: color_data = 12'b111111111111;
20'b01000011010101110111: color_data = 12'b111111111111;
20'b01000011010101111000: color_data = 12'b111111111111;
20'b01000011010101111001: color_data = 12'b111111111111;
20'b01000011010110101101: color_data = 12'b111111111111;
20'b01000011010110101110: color_data = 12'b111111111111;
20'b01000011010110101111: color_data = 12'b111111111111;
20'b01000011010110110000: color_data = 12'b111111111111;
20'b01000011010110110001: color_data = 12'b111111111111;
20'b01000011010110110010: color_data = 12'b111111111111;
20'b01000011010110110011: color_data = 12'b111111111111;
20'b01000011100011110011: color_data = 12'b111111111111;
20'b01000011100011110100: color_data = 12'b111111111111;
20'b01000011100011110101: color_data = 12'b111111111111;
20'b01000011100011110110: color_data = 12'b111111111111;
20'b01000011100011110111: color_data = 12'b111111111111;
20'b01000011100011111000: color_data = 12'b111111111111;
20'b01000011100011111001: color_data = 12'b111111111111;
20'b01000011100011111010: color_data = 12'b111111111111;
20'b01000011100100010101: color_data = 12'b111111111111;
20'b01000011100100010110: color_data = 12'b111111111111;
20'b01000011100100010111: color_data = 12'b111111111111;
20'b01000011100100011000: color_data = 12'b111111111111;
20'b01000011100100011001: color_data = 12'b111111111111;
20'b01000011100100011010: color_data = 12'b111111111111;
20'b01000011100100110100: color_data = 12'b111111111111;
20'b01000011100100110101: color_data = 12'b111111111111;
20'b01000011100100110110: color_data = 12'b111111111111;
20'b01000011100100110111: color_data = 12'b111111111111;
20'b01000011100100111000: color_data = 12'b111111111111;
20'b01000011100100111001: color_data = 12'b111111111111;
20'b01000011100100111010: color_data = 12'b111111111111;
20'b01000011100101001000: color_data = 12'b111111111111;
20'b01000011100101001001: color_data = 12'b111111111111;
20'b01000011100101001010: color_data = 12'b111111111111;
20'b01000011100101001011: color_data = 12'b111111111111;
20'b01000011100101001100: color_data = 12'b111111111111;
20'b01000011100101001101: color_data = 12'b111111111111;
20'b01000011100101010100: color_data = 12'b111111111111;
20'b01000011100101010101: color_data = 12'b111111111111;
20'b01000011100101010110: color_data = 12'b111111111111;
20'b01000011100101010111: color_data = 12'b111111111111;
20'b01000011100101011000: color_data = 12'b111111111111;
20'b01000011100101011001: color_data = 12'b111111111111;
20'b01000011100101011010: color_data = 12'b111111111111;
20'b01000011100101110100: color_data = 12'b111111111111;
20'b01000011100101110101: color_data = 12'b111111111111;
20'b01000011100101110110: color_data = 12'b111111111111;
20'b01000011100101110111: color_data = 12'b111111111111;
20'b01000011100101111000: color_data = 12'b111111111111;
20'b01000011100101111001: color_data = 12'b111111111111;
20'b01000011100110101101: color_data = 12'b111111111111;
20'b01000011100110101110: color_data = 12'b111111111111;
20'b01000011100110101111: color_data = 12'b111111111111;
20'b01000011100110110000: color_data = 12'b111111111111;
20'b01000011100110110001: color_data = 12'b111111111111;
20'b01000011100110110010: color_data = 12'b111111111111;
20'b01000011100110110011: color_data = 12'b111111111111;
20'b01000011110011110011: color_data = 12'b111111111111;
20'b01000011110011110100: color_data = 12'b111111111111;
20'b01000011110011110101: color_data = 12'b111111111111;
20'b01000011110011110110: color_data = 12'b111111111111;
20'b01000011110011110111: color_data = 12'b111111111111;
20'b01000011110011111000: color_data = 12'b111111111111;
20'b01000011110011111001: color_data = 12'b111111111111;
20'b01000011110011111010: color_data = 12'b111111111111;
20'b01000011110100010101: color_data = 12'b111111111111;
20'b01000011110100010110: color_data = 12'b111111111111;
20'b01000011110100010111: color_data = 12'b111111111111;
20'b01000011110100011000: color_data = 12'b111111111111;
20'b01000011110100011001: color_data = 12'b111111111111;
20'b01000011110100011010: color_data = 12'b111111111111;
20'b01000011110100110100: color_data = 12'b111111111111;
20'b01000011110100110101: color_data = 12'b111111111111;
20'b01000011110100110110: color_data = 12'b111111111111;
20'b01000011110100110111: color_data = 12'b111111111111;
20'b01000011110100111000: color_data = 12'b111111111111;
20'b01000011110100111001: color_data = 12'b111111111111;
20'b01000011110100111010: color_data = 12'b111111111111;
20'b01000011110101001000: color_data = 12'b111111111111;
20'b01000011110101001001: color_data = 12'b111111111111;
20'b01000011110101001010: color_data = 12'b111111111111;
20'b01000011110101001011: color_data = 12'b111111111111;
20'b01000011110101001100: color_data = 12'b111111111111;
20'b01000011110101001101: color_data = 12'b111111111111;
20'b01000011110101010100: color_data = 12'b111111111111;
20'b01000011110101010101: color_data = 12'b111111111111;
20'b01000011110101010110: color_data = 12'b111111111111;
20'b01000011110101010111: color_data = 12'b111111111111;
20'b01000011110101011000: color_data = 12'b111111111111;
20'b01000011110101011001: color_data = 12'b111111111111;
20'b01000011110101011010: color_data = 12'b111111111111;
20'b01000011110101110100: color_data = 12'b111111111111;
20'b01000011110101110101: color_data = 12'b111111111111;
20'b01000011110101110110: color_data = 12'b111111111111;
20'b01000011110101110111: color_data = 12'b111111111111;
20'b01000011110101111000: color_data = 12'b111111111111;
20'b01000011110101111001: color_data = 12'b111111111111;
20'b01000011110110101101: color_data = 12'b111111111111;
20'b01000011110110101110: color_data = 12'b111111111111;
20'b01000011110110101111: color_data = 12'b111111111111;
20'b01000011110110110000: color_data = 12'b111111111111;
20'b01000011110110110001: color_data = 12'b111111111111;
20'b01000011110110110010: color_data = 12'b111111111111;
20'b01000011110110110011: color_data = 12'b111111111111;
20'b01000100000011110011: color_data = 12'b111111111111;
20'b01000100000011110100: color_data = 12'b111111111111;
20'b01000100000011110101: color_data = 12'b111111111111;
20'b01000100000011110110: color_data = 12'b111111111111;
20'b01000100000011110111: color_data = 12'b111111111111;
20'b01000100000011111000: color_data = 12'b111111111111;
20'b01000100000011111001: color_data = 12'b111111111111;
20'b01000100000011111010: color_data = 12'b111111111111;
20'b01000100000100010101: color_data = 12'b111111111111;
20'b01000100000100010110: color_data = 12'b111111111111;
20'b01000100000100010111: color_data = 12'b111111111111;
20'b01000100000100011000: color_data = 12'b111111111111;
20'b01000100000100011001: color_data = 12'b111111111111;
20'b01000100000100011010: color_data = 12'b111111111111;
20'b01000100000100110100: color_data = 12'b111111111111;
20'b01000100000100110101: color_data = 12'b111111111111;
20'b01000100000100110110: color_data = 12'b111111111111;
20'b01000100000100110111: color_data = 12'b111111111111;
20'b01000100000100111000: color_data = 12'b111111111111;
20'b01000100000100111001: color_data = 12'b111111111111;
20'b01000100000100111010: color_data = 12'b111111111111;
20'b01000100000101001000: color_data = 12'b111111111111;
20'b01000100000101001001: color_data = 12'b111111111111;
20'b01000100000101001010: color_data = 12'b111111111111;
20'b01000100000101001011: color_data = 12'b111111111111;
20'b01000100000101001100: color_data = 12'b111111111111;
20'b01000100000101001101: color_data = 12'b111111111111;
20'b01000100000101010100: color_data = 12'b111111111111;
20'b01000100000101010101: color_data = 12'b111111111111;
20'b01000100000101010110: color_data = 12'b111111111111;
20'b01000100000101010111: color_data = 12'b111111111111;
20'b01000100000101011000: color_data = 12'b111111111111;
20'b01000100000101011001: color_data = 12'b111111111111;
20'b01000100000101011010: color_data = 12'b111111111111;
20'b01000100000101110100: color_data = 12'b111111111111;
20'b01000100000101110101: color_data = 12'b111111111111;
20'b01000100000101110110: color_data = 12'b111111111111;
20'b01000100000101110111: color_data = 12'b111111111111;
20'b01000100000101111000: color_data = 12'b111111111111;
20'b01000100000101111001: color_data = 12'b111111111111;
20'b01000100000110101101: color_data = 12'b111111111111;
20'b01000100000110101110: color_data = 12'b111111111111;
20'b01000100000110101111: color_data = 12'b111111111111;
20'b01000100000110110000: color_data = 12'b111111111111;
20'b01000100000110110001: color_data = 12'b111111111111;
20'b01000100000110110010: color_data = 12'b111111111111;
20'b01000100000110110011: color_data = 12'b111111111111;
20'b01000100010011011111: color_data = 12'b111111111111;
20'b01000100010011100000: color_data = 12'b111111111111;
20'b01000100010011100001: color_data = 12'b111111111111;
20'b01000100010011100010: color_data = 12'b111111111111;
20'b01000100010011100011: color_data = 12'b111111111111;
20'b01000100010011100100: color_data = 12'b111111111111;
20'b01000100010011100101: color_data = 12'b111111111111;
20'b01000100010011100110: color_data = 12'b111111111111;
20'b01000100010011100111: color_data = 12'b111111111111;
20'b01000100010011101000: color_data = 12'b111111111111;
20'b01000100010011101001: color_data = 12'b111111111111;
20'b01000100010011110011: color_data = 12'b111111111111;
20'b01000100010011110100: color_data = 12'b111111111111;
20'b01000100010011110101: color_data = 12'b111111111111;
20'b01000100010011110110: color_data = 12'b111111111111;
20'b01000100010011110111: color_data = 12'b111111111111;
20'b01000100010011111000: color_data = 12'b111111111111;
20'b01000100010011111001: color_data = 12'b111111111111;
20'b01000100010011111010: color_data = 12'b111111111111;
20'b01000100010100010101: color_data = 12'b111111111111;
20'b01000100010100010110: color_data = 12'b111111111111;
20'b01000100010100010111: color_data = 12'b111111111111;
20'b01000100010100011000: color_data = 12'b111111111111;
20'b01000100010100011001: color_data = 12'b111111111111;
20'b01000100010100011010: color_data = 12'b111111111111;
20'b01000100010100110100: color_data = 12'b111111111111;
20'b01000100010100110101: color_data = 12'b111111111111;
20'b01000100010100110110: color_data = 12'b111111111111;
20'b01000100010100110111: color_data = 12'b111111111111;
20'b01000100010100111000: color_data = 12'b111111111111;
20'b01000100010100111001: color_data = 12'b111111111111;
20'b01000100010100111010: color_data = 12'b111111111111;
20'b01000100010101001000: color_data = 12'b111111111111;
20'b01000100010101001001: color_data = 12'b111111111111;
20'b01000100010101001010: color_data = 12'b111111111111;
20'b01000100010101001011: color_data = 12'b111111111111;
20'b01000100010101001100: color_data = 12'b111111111111;
20'b01000100010101001101: color_data = 12'b111111111111;
20'b01000100010101010100: color_data = 12'b111111111111;
20'b01000100010101010101: color_data = 12'b111111111111;
20'b01000100010101010110: color_data = 12'b111111111111;
20'b01000100010101010111: color_data = 12'b111111111111;
20'b01000100010101011000: color_data = 12'b111111111111;
20'b01000100010101011001: color_data = 12'b111111111111;
20'b01000100010101011010: color_data = 12'b111111111111;
20'b01000100010101110100: color_data = 12'b111111111111;
20'b01000100010101110101: color_data = 12'b111111111111;
20'b01000100010101110110: color_data = 12'b111111111111;
20'b01000100010101110111: color_data = 12'b111111111111;
20'b01000100010101111000: color_data = 12'b111111111111;
20'b01000100010101111001: color_data = 12'b111111111111;
20'b01000100010110101101: color_data = 12'b111111111111;
20'b01000100010110101110: color_data = 12'b111111111111;
20'b01000100010110101111: color_data = 12'b111111111111;
20'b01000100010110110000: color_data = 12'b111111111111;
20'b01000100010110110001: color_data = 12'b111111111111;
20'b01000100010110110010: color_data = 12'b111111111111;
20'b01000100010110110011: color_data = 12'b111111111111;
20'b01000100100011011111: color_data = 12'b111111111111;
20'b01000100100011100000: color_data = 12'b111111111111;
20'b01000100100011100001: color_data = 12'b111111111111;
20'b01000100100011100010: color_data = 12'b111111111111;
20'b01000100100011100011: color_data = 12'b111111111111;
20'b01000100100011100100: color_data = 12'b111111111111;
20'b01000100100011100101: color_data = 12'b111111111111;
20'b01000100100011100110: color_data = 12'b111111111111;
20'b01000100100011100111: color_data = 12'b111111111111;
20'b01000100100011101000: color_data = 12'b111111111111;
20'b01000100100011101001: color_data = 12'b111111111111;
20'b01000100100011110011: color_data = 12'b111111111111;
20'b01000100100011110100: color_data = 12'b111111111111;
20'b01000100100011110101: color_data = 12'b111111111111;
20'b01000100100011110110: color_data = 12'b111111111111;
20'b01000100100011110111: color_data = 12'b111111111111;
20'b01000100100011111000: color_data = 12'b111111111111;
20'b01000100100011111001: color_data = 12'b111111111111;
20'b01000100100011111010: color_data = 12'b111111111111;
20'b01000100100100010101: color_data = 12'b111111111111;
20'b01000100100100010110: color_data = 12'b111111111111;
20'b01000100100100010111: color_data = 12'b111111111111;
20'b01000100100100011000: color_data = 12'b111111111111;
20'b01000100100100011001: color_data = 12'b111111111111;
20'b01000100100100011010: color_data = 12'b111111111111;
20'b01000100100100110100: color_data = 12'b111111111111;
20'b01000100100100110101: color_data = 12'b111111111111;
20'b01000100100100110110: color_data = 12'b111111111111;
20'b01000100100100110111: color_data = 12'b111111111111;
20'b01000100100100111000: color_data = 12'b111111111111;
20'b01000100100100111001: color_data = 12'b111111111111;
20'b01000100100100111010: color_data = 12'b111111111111;
20'b01000100100101001000: color_data = 12'b111111111111;
20'b01000100100101001001: color_data = 12'b111111111111;
20'b01000100100101001010: color_data = 12'b111111111111;
20'b01000100100101001011: color_data = 12'b111111111111;
20'b01000100100101001100: color_data = 12'b111111111111;
20'b01000100100101001101: color_data = 12'b111111111111;
20'b01000100100101010100: color_data = 12'b111111111111;
20'b01000100100101010101: color_data = 12'b111111111111;
20'b01000100100101010110: color_data = 12'b111111111111;
20'b01000100100101010111: color_data = 12'b111111111111;
20'b01000100100101011000: color_data = 12'b111111111111;
20'b01000100100101011001: color_data = 12'b111111111111;
20'b01000100100101011010: color_data = 12'b111111111111;
20'b01000100100101110100: color_data = 12'b111111111111;
20'b01000100100101110101: color_data = 12'b111111111111;
20'b01000100100101110110: color_data = 12'b111111111111;
20'b01000100100101110111: color_data = 12'b111111111111;
20'b01000100100101111000: color_data = 12'b111111111111;
20'b01000100100101111001: color_data = 12'b111111111111;
20'b01000100100110101101: color_data = 12'b111111111111;
20'b01000100100110101110: color_data = 12'b111111111111;
20'b01000100100110101111: color_data = 12'b111111111111;
20'b01000100100110110000: color_data = 12'b111111111111;
20'b01000100100110110001: color_data = 12'b111111111111;
20'b01000100100110110010: color_data = 12'b111111111111;
20'b01000100100110110011: color_data = 12'b111111111111;
20'b01000100110011011111: color_data = 12'b111111111111;
20'b01000100110011100000: color_data = 12'b111111111111;
20'b01000100110011100001: color_data = 12'b111111111111;
20'b01000100110011100010: color_data = 12'b111111111111;
20'b01000100110011100011: color_data = 12'b111111111111;
20'b01000100110011100100: color_data = 12'b111111111111;
20'b01000100110011100101: color_data = 12'b111111111111;
20'b01000100110011100110: color_data = 12'b111111111111;
20'b01000100110011100111: color_data = 12'b111111111111;
20'b01000100110011101000: color_data = 12'b111111111111;
20'b01000100110011101001: color_data = 12'b111111111111;
20'b01000100110011110011: color_data = 12'b111111111111;
20'b01000100110011110100: color_data = 12'b111111111111;
20'b01000100110011110101: color_data = 12'b111111111111;
20'b01000100110011110110: color_data = 12'b111111111111;
20'b01000100110011110111: color_data = 12'b111111111111;
20'b01000100110011111000: color_data = 12'b111111111111;
20'b01000100110011111001: color_data = 12'b111111111111;
20'b01000100110011111010: color_data = 12'b111111111111;
20'b01000100110100010101: color_data = 12'b111111111111;
20'b01000100110100010110: color_data = 12'b111111111111;
20'b01000100110100010111: color_data = 12'b111111111111;
20'b01000100110100011000: color_data = 12'b111111111111;
20'b01000100110100011001: color_data = 12'b111111111111;
20'b01000100110100011010: color_data = 12'b111111111111;
20'b01000100110100011011: color_data = 12'b111111111111;
20'b01000100110100011100: color_data = 12'b111111111111;
20'b01000100110100011101: color_data = 12'b111111111111;
20'b01000100110100011110: color_data = 12'b111111111111;
20'b01000100110100011111: color_data = 12'b111111111111;
20'b01000100110100100000: color_data = 12'b111111111111;
20'b01000100110100100001: color_data = 12'b111111111111;
20'b01000100110100100010: color_data = 12'b111111111111;
20'b01000100110100100011: color_data = 12'b111111111111;
20'b01000100110100100100: color_data = 12'b111111111111;
20'b01000100110100100101: color_data = 12'b111111111111;
20'b01000100110100100110: color_data = 12'b111111111111;
20'b01000100110100100111: color_data = 12'b111111111111;
20'b01000100110100101000: color_data = 12'b111111111111;
20'b01000100110100101001: color_data = 12'b111111111111;
20'b01000100110100101010: color_data = 12'b111111111111;
20'b01000100110100101011: color_data = 12'b111111111111;
20'b01000100110100101100: color_data = 12'b111111111111;
20'b01000100110100101101: color_data = 12'b111111111111;
20'b01000100110100110100: color_data = 12'b111111111111;
20'b01000100110100110101: color_data = 12'b111111111111;
20'b01000100110100110110: color_data = 12'b111111111111;
20'b01000100110100110111: color_data = 12'b111111111111;
20'b01000100110100111000: color_data = 12'b111111111111;
20'b01000100110100111001: color_data = 12'b111111111111;
20'b01000100110100111010: color_data = 12'b111111111111;
20'b01000100110101001000: color_data = 12'b111111111111;
20'b01000100110101001001: color_data = 12'b111111111111;
20'b01000100110101001010: color_data = 12'b111111111111;
20'b01000100110101001011: color_data = 12'b111111111111;
20'b01000100110101001100: color_data = 12'b111111111111;
20'b01000100110101001101: color_data = 12'b111111111111;
20'b01000100110101010100: color_data = 12'b111111111111;
20'b01000100110101010101: color_data = 12'b111111111111;
20'b01000100110101010110: color_data = 12'b111111111111;
20'b01000100110101010111: color_data = 12'b111111111111;
20'b01000100110101011000: color_data = 12'b111111111111;
20'b01000100110101011001: color_data = 12'b111111111111;
20'b01000100110101011010: color_data = 12'b111111111111;
20'b01000100110101011011: color_data = 12'b111111111111;
20'b01000100110101011100: color_data = 12'b111111111111;
20'b01000100110101011101: color_data = 12'b111111111111;
20'b01000100110101011110: color_data = 12'b111111111111;
20'b01000100110101011111: color_data = 12'b111111111111;
20'b01000100110101100000: color_data = 12'b111111111111;
20'b01000100110101100001: color_data = 12'b111111111111;
20'b01000100110101100010: color_data = 12'b111111111111;
20'b01000100110101100011: color_data = 12'b111111111111;
20'b01000100110101100100: color_data = 12'b111111111111;
20'b01000100110101100101: color_data = 12'b111111111111;
20'b01000100110101100110: color_data = 12'b111111111111;
20'b01000100110101100111: color_data = 12'b111111111111;
20'b01000100110101101000: color_data = 12'b111111111111;
20'b01000100110101101001: color_data = 12'b111111111111;
20'b01000100110101101010: color_data = 12'b111111111111;
20'b01000100110101101011: color_data = 12'b111111111111;
20'b01000100110101101100: color_data = 12'b111111111111;
20'b01000100110101101101: color_data = 12'b111111111111;
20'b01000100110101110100: color_data = 12'b111111111111;
20'b01000100110101110101: color_data = 12'b111111111111;
20'b01000100110101110110: color_data = 12'b111111111111;
20'b01000100110101110111: color_data = 12'b111111111111;
20'b01000100110101111000: color_data = 12'b111111111111;
20'b01000100110101111001: color_data = 12'b111111111111;
20'b01000100110110011010: color_data = 12'b111111111111;
20'b01000100110110011011: color_data = 12'b111111111111;
20'b01000100110110011100: color_data = 12'b111111111111;
20'b01000100110110011101: color_data = 12'b111111111111;
20'b01000100110110011110: color_data = 12'b111111111111;
20'b01000100110110011111: color_data = 12'b111111111111;
20'b01000100110110100000: color_data = 12'b111111111111;
20'b01000100110110100001: color_data = 12'b111111111111;
20'b01000100110110100010: color_data = 12'b111111111111;
20'b01000100110110100011: color_data = 12'b111111111111;
20'b01000100110110100100: color_data = 12'b111111111111;
20'b01000100110110100101: color_data = 12'b111111111111;
20'b01000100110110100110: color_data = 12'b111111111111;
20'b01000100110110100111: color_data = 12'b111111111111;
20'b01000100110110101000: color_data = 12'b111111111111;
20'b01000100110110101001: color_data = 12'b111111111111;
20'b01000100110110101010: color_data = 12'b111111111111;
20'b01000100110110101011: color_data = 12'b111111111111;
20'b01000100110110101100: color_data = 12'b111111111111;
20'b01000100110110101101: color_data = 12'b111111111111;
20'b01000100110110101110: color_data = 12'b111111111111;
20'b01000100110110101111: color_data = 12'b111111111111;
20'b01000100110110110000: color_data = 12'b111111111111;
20'b01000100110110110001: color_data = 12'b111111111111;
20'b01000100110110110010: color_data = 12'b111111111111;
20'b01000100110110110011: color_data = 12'b111111111111;
20'b01000101000011011111: color_data = 12'b111111111111;
20'b01000101000011100000: color_data = 12'b111111111111;
20'b01000101000011100001: color_data = 12'b111111111111;
20'b01000101000011100010: color_data = 12'b111111111111;
20'b01000101000011100011: color_data = 12'b111111111111;
20'b01000101000011100100: color_data = 12'b111111111111;
20'b01000101000011100101: color_data = 12'b111111111111;
20'b01000101000011100110: color_data = 12'b111111111111;
20'b01000101000011100111: color_data = 12'b111111111111;
20'b01000101000011101000: color_data = 12'b111111111111;
20'b01000101000011101001: color_data = 12'b111111111111;
20'b01000101000011110011: color_data = 12'b111111111111;
20'b01000101000011110100: color_data = 12'b111111111111;
20'b01000101000011110101: color_data = 12'b111111111111;
20'b01000101000011110110: color_data = 12'b111111111111;
20'b01000101000011110111: color_data = 12'b111111111111;
20'b01000101000011111000: color_data = 12'b111111111111;
20'b01000101000011111001: color_data = 12'b111111111111;
20'b01000101000011111010: color_data = 12'b111111111111;
20'b01000101000100010101: color_data = 12'b111111111111;
20'b01000101000100010110: color_data = 12'b111111111111;
20'b01000101000100010111: color_data = 12'b111111111111;
20'b01000101000100011000: color_data = 12'b111111111111;
20'b01000101000100011001: color_data = 12'b111111111111;
20'b01000101000100011010: color_data = 12'b111111111111;
20'b01000101000100011011: color_data = 12'b111111111111;
20'b01000101000100011100: color_data = 12'b111111111111;
20'b01000101000100011101: color_data = 12'b111111111111;
20'b01000101000100011110: color_data = 12'b111111111111;
20'b01000101000100011111: color_data = 12'b111111111111;
20'b01000101000100100000: color_data = 12'b111111111111;
20'b01000101000100100001: color_data = 12'b111111111111;
20'b01000101000100100010: color_data = 12'b111111111111;
20'b01000101000100100011: color_data = 12'b111111111111;
20'b01000101000100100100: color_data = 12'b111111111111;
20'b01000101000100100101: color_data = 12'b111111111111;
20'b01000101000100100110: color_data = 12'b111111111111;
20'b01000101000100100111: color_data = 12'b111111111111;
20'b01000101000100101000: color_data = 12'b111111111111;
20'b01000101000100101001: color_data = 12'b111111111111;
20'b01000101000100101010: color_data = 12'b111111111111;
20'b01000101000100101011: color_data = 12'b111111111111;
20'b01000101000100101100: color_data = 12'b111111111111;
20'b01000101000100101101: color_data = 12'b111111111111;
20'b01000101000100110100: color_data = 12'b111111111111;
20'b01000101000100110101: color_data = 12'b111111111111;
20'b01000101000100110110: color_data = 12'b111111111111;
20'b01000101000100110111: color_data = 12'b111111111111;
20'b01000101000100111000: color_data = 12'b111111111111;
20'b01000101000100111001: color_data = 12'b111111111111;
20'b01000101000100111010: color_data = 12'b111111111111;
20'b01000101000101001000: color_data = 12'b111111111111;
20'b01000101000101001001: color_data = 12'b111111111111;
20'b01000101000101001010: color_data = 12'b111111111111;
20'b01000101000101001011: color_data = 12'b111111111111;
20'b01000101000101001100: color_data = 12'b111111111111;
20'b01000101000101001101: color_data = 12'b111111111111;
20'b01000101000101010100: color_data = 12'b111111111111;
20'b01000101000101010101: color_data = 12'b111111111111;
20'b01000101000101010110: color_data = 12'b111111111111;
20'b01000101000101010111: color_data = 12'b111111111111;
20'b01000101000101011000: color_data = 12'b111111111111;
20'b01000101000101011001: color_data = 12'b111111111111;
20'b01000101000101011010: color_data = 12'b111111111111;
20'b01000101000101011011: color_data = 12'b111111111111;
20'b01000101000101011100: color_data = 12'b111111111111;
20'b01000101000101011101: color_data = 12'b111111111111;
20'b01000101000101011110: color_data = 12'b111111111111;
20'b01000101000101011111: color_data = 12'b111111111111;
20'b01000101000101100000: color_data = 12'b111111111111;
20'b01000101000101100001: color_data = 12'b111111111111;
20'b01000101000101100010: color_data = 12'b111111111111;
20'b01000101000101100011: color_data = 12'b111111111111;
20'b01000101000101100100: color_data = 12'b111111111111;
20'b01000101000101100101: color_data = 12'b111111111111;
20'b01000101000101100110: color_data = 12'b111111111111;
20'b01000101000101100111: color_data = 12'b111111111111;
20'b01000101000101101000: color_data = 12'b111111111111;
20'b01000101000101101001: color_data = 12'b111111111111;
20'b01000101000101101010: color_data = 12'b111111111111;
20'b01000101000101101011: color_data = 12'b111111111111;
20'b01000101000101101100: color_data = 12'b111111111111;
20'b01000101000101101101: color_data = 12'b111111111111;
20'b01000101000101110100: color_data = 12'b111111111111;
20'b01000101000101110101: color_data = 12'b111111111111;
20'b01000101000101110110: color_data = 12'b111111111111;
20'b01000101000101110111: color_data = 12'b111111111111;
20'b01000101000101111000: color_data = 12'b111111111111;
20'b01000101000101111001: color_data = 12'b111111111111;
20'b01000101000110011010: color_data = 12'b111111111111;
20'b01000101000110011011: color_data = 12'b111111111111;
20'b01000101000110011100: color_data = 12'b111111111111;
20'b01000101000110011101: color_data = 12'b111111111111;
20'b01000101000110011110: color_data = 12'b111111111111;
20'b01000101000110011111: color_data = 12'b111111111111;
20'b01000101000110100000: color_data = 12'b111111111111;
20'b01000101000110100001: color_data = 12'b111111111111;
20'b01000101000110100010: color_data = 12'b111111111111;
20'b01000101000110100011: color_data = 12'b111111111111;
20'b01000101000110100100: color_data = 12'b111111111111;
20'b01000101000110100101: color_data = 12'b111111111111;
20'b01000101000110100110: color_data = 12'b111111111111;
20'b01000101000110100111: color_data = 12'b111111111111;
20'b01000101000110101000: color_data = 12'b111111111111;
20'b01000101000110101001: color_data = 12'b111111111111;
20'b01000101000110101010: color_data = 12'b111111111111;
20'b01000101000110101011: color_data = 12'b111111111111;
20'b01000101000110101100: color_data = 12'b111111111111;
20'b01000101000110101101: color_data = 12'b111111111111;
20'b01000101000110101110: color_data = 12'b111111111111;
20'b01000101000110101111: color_data = 12'b111111111111;
20'b01000101000110110000: color_data = 12'b111111111111;
20'b01000101000110110001: color_data = 12'b111111111111;
20'b01000101000110110010: color_data = 12'b111111111111;
20'b01000101000110110011: color_data = 12'b111111111111;
20'b01000101010011011111: color_data = 12'b111111111111;
20'b01000101010011100000: color_data = 12'b111111111111;
20'b01000101010011100001: color_data = 12'b111111111111;
20'b01000101010011100010: color_data = 12'b111111111111;
20'b01000101010011100011: color_data = 12'b111111111111;
20'b01000101010011100100: color_data = 12'b111111111111;
20'b01000101010011100101: color_data = 12'b111111111111;
20'b01000101010011100110: color_data = 12'b111111111111;
20'b01000101010011100111: color_data = 12'b111111111111;
20'b01000101010011101000: color_data = 12'b111111111111;
20'b01000101010011101001: color_data = 12'b111111111111;
20'b01000101010011110011: color_data = 12'b111111111111;
20'b01000101010011110100: color_data = 12'b111111111111;
20'b01000101010011110101: color_data = 12'b111111111111;
20'b01000101010011110110: color_data = 12'b111111111111;
20'b01000101010011110111: color_data = 12'b111111111111;
20'b01000101010011111000: color_data = 12'b111111111111;
20'b01000101010011111001: color_data = 12'b111111111111;
20'b01000101010011111010: color_data = 12'b111111111111;
20'b01000101010100010101: color_data = 12'b111111111111;
20'b01000101010100010110: color_data = 12'b111111111111;
20'b01000101010100010111: color_data = 12'b111111111111;
20'b01000101010100011000: color_data = 12'b111111111111;
20'b01000101010100011001: color_data = 12'b111111111111;
20'b01000101010100011010: color_data = 12'b111111111111;
20'b01000101010100011011: color_data = 12'b111111111111;
20'b01000101010100011100: color_data = 12'b111111111111;
20'b01000101010100011101: color_data = 12'b111111111111;
20'b01000101010100011110: color_data = 12'b111111111111;
20'b01000101010100011111: color_data = 12'b111111111111;
20'b01000101010100100000: color_data = 12'b111111111111;
20'b01000101010100100001: color_data = 12'b111111111111;
20'b01000101010100100010: color_data = 12'b111111111111;
20'b01000101010100100011: color_data = 12'b111111111111;
20'b01000101010100100100: color_data = 12'b111111111111;
20'b01000101010100100101: color_data = 12'b111111111111;
20'b01000101010100100110: color_data = 12'b111111111111;
20'b01000101010100100111: color_data = 12'b111111111111;
20'b01000101010100101000: color_data = 12'b111111111111;
20'b01000101010100101001: color_data = 12'b111111111111;
20'b01000101010100101010: color_data = 12'b111111111111;
20'b01000101010100101011: color_data = 12'b111111111111;
20'b01000101010100101100: color_data = 12'b111111111111;
20'b01000101010100101101: color_data = 12'b111111111111;
20'b01000101010100110100: color_data = 12'b111111111111;
20'b01000101010100110101: color_data = 12'b111111111111;
20'b01000101010100110110: color_data = 12'b111111111111;
20'b01000101010100110111: color_data = 12'b111111111111;
20'b01000101010100111000: color_data = 12'b111111111111;
20'b01000101010100111001: color_data = 12'b111111111111;
20'b01000101010100111010: color_data = 12'b111111111111;
20'b01000101010101001000: color_data = 12'b111111111111;
20'b01000101010101001001: color_data = 12'b111111111111;
20'b01000101010101001010: color_data = 12'b111111111111;
20'b01000101010101001011: color_data = 12'b111111111111;
20'b01000101010101001100: color_data = 12'b111111111111;
20'b01000101010101001101: color_data = 12'b111111111111;
20'b01000101010101010100: color_data = 12'b111111111111;
20'b01000101010101010101: color_data = 12'b111111111111;
20'b01000101010101010110: color_data = 12'b111111111111;
20'b01000101010101010111: color_data = 12'b111111111111;
20'b01000101010101011000: color_data = 12'b111111111111;
20'b01000101010101011001: color_data = 12'b111111111111;
20'b01000101010101011010: color_data = 12'b111111111111;
20'b01000101010101011011: color_data = 12'b111111111111;
20'b01000101010101011100: color_data = 12'b111111111111;
20'b01000101010101011101: color_data = 12'b111111111111;
20'b01000101010101011110: color_data = 12'b111111111111;
20'b01000101010101011111: color_data = 12'b111111111111;
20'b01000101010101100000: color_data = 12'b111111111111;
20'b01000101010101100001: color_data = 12'b111111111111;
20'b01000101010101100010: color_data = 12'b111111111111;
20'b01000101010101100011: color_data = 12'b111111111111;
20'b01000101010101100100: color_data = 12'b111111111111;
20'b01000101010101100101: color_data = 12'b111111111111;
20'b01000101010101100110: color_data = 12'b111111111111;
20'b01000101010101100111: color_data = 12'b111111111111;
20'b01000101010101101000: color_data = 12'b111111111111;
20'b01000101010101101001: color_data = 12'b111111111111;
20'b01000101010101101010: color_data = 12'b111111111111;
20'b01000101010101101011: color_data = 12'b111111111111;
20'b01000101010101101100: color_data = 12'b111111111111;
20'b01000101010101101101: color_data = 12'b111111111111;
20'b01000101010101110100: color_data = 12'b111111111111;
20'b01000101010101110101: color_data = 12'b111111111111;
20'b01000101010101110110: color_data = 12'b111111111111;
20'b01000101010101110111: color_data = 12'b111111111111;
20'b01000101010101111000: color_data = 12'b111111111111;
20'b01000101010101111001: color_data = 12'b111111111111;
20'b01000101010110011010: color_data = 12'b111111111111;
20'b01000101010110011011: color_data = 12'b111111111111;
20'b01000101010110011100: color_data = 12'b111111111111;
20'b01000101010110011101: color_data = 12'b111111111111;
20'b01000101010110011110: color_data = 12'b111111111111;
20'b01000101010110011111: color_data = 12'b111111111111;
20'b01000101010110100000: color_data = 12'b111111111111;
20'b01000101010110100001: color_data = 12'b111111111111;
20'b01000101010110100010: color_data = 12'b111111111111;
20'b01000101010110100011: color_data = 12'b111111111111;
20'b01000101010110100100: color_data = 12'b111111111111;
20'b01000101010110100101: color_data = 12'b111111111111;
20'b01000101010110100110: color_data = 12'b111111111111;
20'b01000101010110100111: color_data = 12'b111111111111;
20'b01000101010110101000: color_data = 12'b111111111111;
20'b01000101010110101001: color_data = 12'b111111111111;
20'b01000101010110101010: color_data = 12'b111111111111;
20'b01000101010110101011: color_data = 12'b111111111111;
20'b01000101010110101100: color_data = 12'b111111111111;
20'b01000101010110101101: color_data = 12'b111111111111;
20'b01000101010110101110: color_data = 12'b111111111111;
20'b01000101010110101111: color_data = 12'b111111111111;
20'b01000101010110110000: color_data = 12'b111111111111;
20'b01000101010110110001: color_data = 12'b111111111111;
20'b01000101010110110010: color_data = 12'b111111111111;
20'b01000101010110110011: color_data = 12'b111111111111;
20'b01000101100011011111: color_data = 12'b111111111111;
20'b01000101100011100000: color_data = 12'b111111111111;
20'b01000101100011100001: color_data = 12'b111111111111;
20'b01000101100011100010: color_data = 12'b111111111111;
20'b01000101100011100011: color_data = 12'b111111111111;
20'b01000101100011100100: color_data = 12'b111111111111;
20'b01000101100011100101: color_data = 12'b111111111111;
20'b01000101100011100110: color_data = 12'b111111111111;
20'b01000101100011100111: color_data = 12'b111111111111;
20'b01000101100011101000: color_data = 12'b111111111111;
20'b01000101100011101001: color_data = 12'b111111111111;
20'b01000101100011110011: color_data = 12'b111111111111;
20'b01000101100011110100: color_data = 12'b111111111111;
20'b01000101100011110101: color_data = 12'b111111111111;
20'b01000101100011110110: color_data = 12'b111111111111;
20'b01000101100011110111: color_data = 12'b111111111111;
20'b01000101100011111000: color_data = 12'b111111111111;
20'b01000101100011111001: color_data = 12'b111111111111;
20'b01000101100011111010: color_data = 12'b111111111111;
20'b01000101100100010101: color_data = 12'b111111111111;
20'b01000101100100010110: color_data = 12'b111111111111;
20'b01000101100100010111: color_data = 12'b111111111111;
20'b01000101100100011000: color_data = 12'b111111111111;
20'b01000101100100011001: color_data = 12'b111111111111;
20'b01000101100100011010: color_data = 12'b111111111111;
20'b01000101100100011011: color_data = 12'b111111111111;
20'b01000101100100011100: color_data = 12'b111111111111;
20'b01000101100100011101: color_data = 12'b111111111111;
20'b01000101100100011110: color_data = 12'b111111111111;
20'b01000101100100011111: color_data = 12'b111111111111;
20'b01000101100100100000: color_data = 12'b111111111111;
20'b01000101100100100001: color_data = 12'b111111111111;
20'b01000101100100100010: color_data = 12'b111111111111;
20'b01000101100100100011: color_data = 12'b111111111111;
20'b01000101100100100100: color_data = 12'b111111111111;
20'b01000101100100100101: color_data = 12'b111111111111;
20'b01000101100100100110: color_data = 12'b111111111111;
20'b01000101100100100111: color_data = 12'b111111111111;
20'b01000101100100101000: color_data = 12'b111111111111;
20'b01000101100100101001: color_data = 12'b111111111111;
20'b01000101100100101010: color_data = 12'b111111111111;
20'b01000101100100101011: color_data = 12'b111111111111;
20'b01000101100100101100: color_data = 12'b111111111111;
20'b01000101100100101101: color_data = 12'b111111111111;
20'b01000101100100110100: color_data = 12'b111111111111;
20'b01000101100100110101: color_data = 12'b111111111111;
20'b01000101100100110110: color_data = 12'b111111111111;
20'b01000101100100110111: color_data = 12'b111111111111;
20'b01000101100100111000: color_data = 12'b111111111111;
20'b01000101100100111001: color_data = 12'b111111111111;
20'b01000101100100111010: color_data = 12'b111111111111;
20'b01000101100101001000: color_data = 12'b111111111111;
20'b01000101100101001001: color_data = 12'b111111111111;
20'b01000101100101001010: color_data = 12'b111111111111;
20'b01000101100101001011: color_data = 12'b111111111111;
20'b01000101100101001100: color_data = 12'b111111111111;
20'b01000101100101001101: color_data = 12'b111111111111;
20'b01000101100101010100: color_data = 12'b111111111111;
20'b01000101100101010101: color_data = 12'b111111111111;
20'b01000101100101010110: color_data = 12'b111111111111;
20'b01000101100101010111: color_data = 12'b111111111111;
20'b01000101100101011000: color_data = 12'b111111111111;
20'b01000101100101011001: color_data = 12'b111111111111;
20'b01000101100101011010: color_data = 12'b111111111111;
20'b01000101100101011011: color_data = 12'b111111111111;
20'b01000101100101011100: color_data = 12'b111111111111;
20'b01000101100101011101: color_data = 12'b111111111111;
20'b01000101100101011110: color_data = 12'b111111111111;
20'b01000101100101011111: color_data = 12'b111111111111;
20'b01000101100101100000: color_data = 12'b111111111111;
20'b01000101100101100001: color_data = 12'b111111111111;
20'b01000101100101100010: color_data = 12'b111111111111;
20'b01000101100101100011: color_data = 12'b111111111111;
20'b01000101100101100100: color_data = 12'b111111111111;
20'b01000101100101100101: color_data = 12'b111111111111;
20'b01000101100101100110: color_data = 12'b111111111111;
20'b01000101100101100111: color_data = 12'b111111111111;
20'b01000101100101101000: color_data = 12'b111111111111;
20'b01000101100101101001: color_data = 12'b111111111111;
20'b01000101100101101010: color_data = 12'b111111111111;
20'b01000101100101101011: color_data = 12'b111111111111;
20'b01000101100101101100: color_data = 12'b111111111111;
20'b01000101100101101101: color_data = 12'b111111111111;
20'b01000101100101110100: color_data = 12'b111111111111;
20'b01000101100101110101: color_data = 12'b111111111111;
20'b01000101100101110110: color_data = 12'b111111111111;
20'b01000101100101110111: color_data = 12'b111111111111;
20'b01000101100101111000: color_data = 12'b111111111111;
20'b01000101100101111001: color_data = 12'b111111111111;
20'b01000101100110011010: color_data = 12'b111111111111;
20'b01000101100110011011: color_data = 12'b111111111111;
20'b01000101100110011100: color_data = 12'b111111111111;
20'b01000101100110011101: color_data = 12'b111111111111;
20'b01000101100110011110: color_data = 12'b111111111111;
20'b01000101100110011111: color_data = 12'b111111111111;
20'b01000101100110100000: color_data = 12'b111111111111;
20'b01000101100110100001: color_data = 12'b111111111111;
20'b01000101100110100010: color_data = 12'b111111111111;
20'b01000101100110100011: color_data = 12'b111111111111;
20'b01000101100110100100: color_data = 12'b111111111111;
20'b01000101100110100101: color_data = 12'b111111111111;
20'b01000101100110100110: color_data = 12'b111111111111;
20'b01000101100110100111: color_data = 12'b111111111111;
20'b01000101100110101000: color_data = 12'b111111111111;
20'b01000101100110101001: color_data = 12'b111111111111;
20'b01000101100110101010: color_data = 12'b111111111111;
20'b01000101100110101011: color_data = 12'b111111111111;
20'b01000101100110101100: color_data = 12'b111111111111;
20'b01000101100110101101: color_data = 12'b111111111111;
20'b01000101100110101110: color_data = 12'b111111111111;
20'b01000101100110101111: color_data = 12'b111111111111;
20'b01000101100110110000: color_data = 12'b111111111111;
20'b01000101100110110001: color_data = 12'b111111111111;
20'b01000101100110110010: color_data = 12'b111111111111;
20'b01000101100110110011: color_data = 12'b111111111111;
20'b01000101110011011111: color_data = 12'b111111111111;
20'b01000101110011100000: color_data = 12'b111111111111;
20'b01000101110011100001: color_data = 12'b111111111111;
20'b01000101110011100010: color_data = 12'b111111111111;
20'b01000101110011100011: color_data = 12'b111111111111;
20'b01000101110011100100: color_data = 12'b111111111111;
20'b01000101110011100101: color_data = 12'b111111111111;
20'b01000101110011100110: color_data = 12'b111111111111;
20'b01000101110011100111: color_data = 12'b111111111111;
20'b01000101110011101000: color_data = 12'b111111111111;
20'b01000101110011101001: color_data = 12'b111111111111;
20'b01000101110011110011: color_data = 12'b111111111111;
20'b01000101110011110100: color_data = 12'b111111111111;
20'b01000101110011110101: color_data = 12'b111111111111;
20'b01000101110011110110: color_data = 12'b111111111111;
20'b01000101110011110111: color_data = 12'b111111111111;
20'b01000101110011111000: color_data = 12'b111111111111;
20'b01000101110011111001: color_data = 12'b111111111111;
20'b01000101110011111010: color_data = 12'b111111111111;
20'b01000101110100010101: color_data = 12'b111111111111;
20'b01000101110100010110: color_data = 12'b111111111111;
20'b01000101110100010111: color_data = 12'b111111111111;
20'b01000101110100011000: color_data = 12'b111111111111;
20'b01000101110100011001: color_data = 12'b111111111111;
20'b01000101110100011010: color_data = 12'b111111111111;
20'b01000101110100011011: color_data = 12'b111111111111;
20'b01000101110100011100: color_data = 12'b111111111111;
20'b01000101110100011101: color_data = 12'b111111111111;
20'b01000101110100011110: color_data = 12'b111111111111;
20'b01000101110100011111: color_data = 12'b111111111111;
20'b01000101110100100000: color_data = 12'b111111111111;
20'b01000101110100100001: color_data = 12'b111111111111;
20'b01000101110100100010: color_data = 12'b111111111111;
20'b01000101110100100011: color_data = 12'b111111111111;
20'b01000101110100100100: color_data = 12'b111111111111;
20'b01000101110100100101: color_data = 12'b111111111111;
20'b01000101110100100110: color_data = 12'b111111111111;
20'b01000101110100100111: color_data = 12'b111111111111;
20'b01000101110100101000: color_data = 12'b111111111111;
20'b01000101110100101001: color_data = 12'b111111111111;
20'b01000101110100101010: color_data = 12'b111111111111;
20'b01000101110100101011: color_data = 12'b111111111111;
20'b01000101110100101100: color_data = 12'b111111111111;
20'b01000101110100101101: color_data = 12'b111111111111;
20'b01000101110100110100: color_data = 12'b111111111111;
20'b01000101110100110101: color_data = 12'b111111111111;
20'b01000101110100110110: color_data = 12'b111111111111;
20'b01000101110100110111: color_data = 12'b111111111111;
20'b01000101110100111000: color_data = 12'b111111111111;
20'b01000101110100111001: color_data = 12'b111111111111;
20'b01000101110100111010: color_data = 12'b111111111111;
20'b01000101110101001000: color_data = 12'b111111111111;
20'b01000101110101001001: color_data = 12'b111111111111;
20'b01000101110101001010: color_data = 12'b111111111111;
20'b01000101110101001011: color_data = 12'b111111111111;
20'b01000101110101001100: color_data = 12'b111111111111;
20'b01000101110101001101: color_data = 12'b111111111111;
20'b01000101110101010100: color_data = 12'b111111111111;
20'b01000101110101010101: color_data = 12'b111111111111;
20'b01000101110101010110: color_data = 12'b111111111111;
20'b01000101110101010111: color_data = 12'b111111111111;
20'b01000101110101011000: color_data = 12'b111111111111;
20'b01000101110101011001: color_data = 12'b111111111111;
20'b01000101110101011010: color_data = 12'b111111111111;
20'b01000101110101011011: color_data = 12'b111111111111;
20'b01000101110101011100: color_data = 12'b111111111111;
20'b01000101110101011101: color_data = 12'b111111111111;
20'b01000101110101011110: color_data = 12'b111111111111;
20'b01000101110101011111: color_data = 12'b111111111111;
20'b01000101110101100000: color_data = 12'b111111111111;
20'b01000101110101100001: color_data = 12'b111111111111;
20'b01000101110101100010: color_data = 12'b111111111111;
20'b01000101110101100011: color_data = 12'b111111111111;
20'b01000101110101100100: color_data = 12'b111111111111;
20'b01000101110101100101: color_data = 12'b111111111111;
20'b01000101110101100110: color_data = 12'b111111111111;
20'b01000101110101100111: color_data = 12'b111111111111;
20'b01000101110101101000: color_data = 12'b111111111111;
20'b01000101110101101001: color_data = 12'b111111111111;
20'b01000101110101101010: color_data = 12'b111111111111;
20'b01000101110101101011: color_data = 12'b111111111111;
20'b01000101110101101100: color_data = 12'b111111111111;
20'b01000101110101101101: color_data = 12'b111111111111;
20'b01000101110101110100: color_data = 12'b111111111111;
20'b01000101110101110101: color_data = 12'b111111111111;
20'b01000101110101110110: color_data = 12'b111111111111;
20'b01000101110101110111: color_data = 12'b111111111111;
20'b01000101110101111000: color_data = 12'b111111111111;
20'b01000101110101111001: color_data = 12'b111111111111;
20'b01000101110110011010: color_data = 12'b111111111111;
20'b01000101110110011011: color_data = 12'b111111111111;
20'b01000101110110011100: color_data = 12'b111111111111;
20'b01000101110110011101: color_data = 12'b111111111111;
20'b01000101110110011110: color_data = 12'b111111111111;
20'b01000101110110011111: color_data = 12'b111111111111;
20'b01000101110110100000: color_data = 12'b111111111111;
20'b01000101110110100001: color_data = 12'b111111111111;
20'b01000101110110100010: color_data = 12'b111111111111;
20'b01000101110110100011: color_data = 12'b111111111111;
20'b01000101110110100100: color_data = 12'b111111111111;
20'b01000101110110100101: color_data = 12'b111111111111;
20'b01000101110110100110: color_data = 12'b111111111111;
20'b01000101110110100111: color_data = 12'b111111111111;
20'b01000101110110101000: color_data = 12'b111111111111;
20'b01000101110110101001: color_data = 12'b111111111111;
20'b01000101110110101010: color_data = 12'b111111111111;
20'b01000101110110101011: color_data = 12'b111111111111;
20'b01000101110110101100: color_data = 12'b111111111111;
20'b01000101110110101101: color_data = 12'b111111111111;
20'b01000101110110101110: color_data = 12'b111111111111;
20'b01000101110110101111: color_data = 12'b111111111111;
20'b01000101110110110000: color_data = 12'b111111111111;
20'b01000101110110110001: color_data = 12'b111111111111;
20'b01000101110110110010: color_data = 12'b111111111111;
20'b01000101110110110011: color_data = 12'b111111111111;
20'b01000110000011011111: color_data = 12'b111111111111;
20'b01000110000011100000: color_data = 12'b111111111111;
20'b01000110000011100001: color_data = 12'b111111111111;
20'b01000110000011100010: color_data = 12'b111111111111;
20'b01000110000011100011: color_data = 12'b111111111111;
20'b01000110000011100100: color_data = 12'b111111111111;
20'b01000110000011100101: color_data = 12'b111111111111;
20'b01000110000011100110: color_data = 12'b111111111111;
20'b01000110000011100111: color_data = 12'b111111111111;
20'b01000110000011101000: color_data = 12'b111111111111;
20'b01000110000011101001: color_data = 12'b111111111111;
20'b01000110000011110011: color_data = 12'b111111111111;
20'b01000110000011110100: color_data = 12'b111111111111;
20'b01000110000011110101: color_data = 12'b111111111111;
20'b01000110000011110110: color_data = 12'b111111111111;
20'b01000110000011110111: color_data = 12'b111111111111;
20'b01000110000011111000: color_data = 12'b111111111111;
20'b01000110000011111001: color_data = 12'b111111111111;
20'b01000110000011111010: color_data = 12'b111111111111;
20'b01000110000100010101: color_data = 12'b111111111111;
20'b01000110000100010110: color_data = 12'b111111111111;
20'b01000110000100010111: color_data = 12'b111111111111;
20'b01000110000100011000: color_data = 12'b111111111111;
20'b01000110000100011001: color_data = 12'b111111111111;
20'b01000110000100011010: color_data = 12'b111111111111;
20'b01000110000100011011: color_data = 12'b111111111111;
20'b01000110000100011100: color_data = 12'b111111111111;
20'b01000110000100011101: color_data = 12'b111111111111;
20'b01000110000100011110: color_data = 12'b111111111111;
20'b01000110000100011111: color_data = 12'b111111111111;
20'b01000110000100100000: color_data = 12'b111111111111;
20'b01000110000100100001: color_data = 12'b111111111111;
20'b01000110000100100010: color_data = 12'b111111111111;
20'b01000110000100100011: color_data = 12'b111111111111;
20'b01000110000100100100: color_data = 12'b111111111111;
20'b01000110000100100101: color_data = 12'b111111111111;
20'b01000110000100100110: color_data = 12'b111111111111;
20'b01000110000100100111: color_data = 12'b111111111111;
20'b01000110000100101000: color_data = 12'b111111111111;
20'b01000110000100101001: color_data = 12'b111111111111;
20'b01000110000100101010: color_data = 12'b111111111111;
20'b01000110000100101011: color_data = 12'b111111111111;
20'b01000110000100101100: color_data = 12'b111111111111;
20'b01000110000100101101: color_data = 12'b111111111111;
20'b01000110000100110100: color_data = 12'b111111111111;
20'b01000110000100110101: color_data = 12'b111111111111;
20'b01000110000100110110: color_data = 12'b111111111111;
20'b01000110000100110111: color_data = 12'b111111111111;
20'b01000110000100111000: color_data = 12'b111111111111;
20'b01000110000100111001: color_data = 12'b111111111111;
20'b01000110000100111010: color_data = 12'b111111111111;
20'b01000110000101001000: color_data = 12'b111111111111;
20'b01000110000101001001: color_data = 12'b111111111111;
20'b01000110000101001010: color_data = 12'b111111111111;
20'b01000110000101001011: color_data = 12'b111111111111;
20'b01000110000101001100: color_data = 12'b111111111111;
20'b01000110000101001101: color_data = 12'b111111111111;
20'b01000110000101010100: color_data = 12'b111111111111;
20'b01000110000101010101: color_data = 12'b111111111111;
20'b01000110000101010110: color_data = 12'b111111111111;
20'b01000110000101010111: color_data = 12'b111111111111;
20'b01000110000101011000: color_data = 12'b111111111111;
20'b01000110000101011001: color_data = 12'b111111111111;
20'b01000110000101011010: color_data = 12'b111111111111;
20'b01000110000101011011: color_data = 12'b111111111111;
20'b01000110000101011100: color_data = 12'b111111111111;
20'b01000110000101011101: color_data = 12'b111111111111;
20'b01000110000101011110: color_data = 12'b111111111111;
20'b01000110000101011111: color_data = 12'b111111111111;
20'b01000110000101100000: color_data = 12'b111111111111;
20'b01000110000101100001: color_data = 12'b111111111111;
20'b01000110000101100010: color_data = 12'b111111111111;
20'b01000110000101100011: color_data = 12'b111111111111;
20'b01000110000101100100: color_data = 12'b111111111111;
20'b01000110000101100101: color_data = 12'b111111111111;
20'b01000110000101100110: color_data = 12'b111111111111;
20'b01000110000101100111: color_data = 12'b111111111111;
20'b01000110000101101000: color_data = 12'b111111111111;
20'b01000110000101101001: color_data = 12'b111111111111;
20'b01000110000101101010: color_data = 12'b111111111111;
20'b01000110000101101011: color_data = 12'b111111111111;
20'b01000110000101101100: color_data = 12'b111111111111;
20'b01000110000101101101: color_data = 12'b111111111111;
20'b01000110000101110100: color_data = 12'b111111111111;
20'b01000110000101110101: color_data = 12'b111111111111;
20'b01000110000101110110: color_data = 12'b111111111111;
20'b01000110000101110111: color_data = 12'b111111111111;
20'b01000110000101111000: color_data = 12'b111111111111;
20'b01000110000101111001: color_data = 12'b111111111111;
20'b01000110000110011010: color_data = 12'b111111111111;
20'b01000110000110011011: color_data = 12'b111111111111;
20'b01000110000110011100: color_data = 12'b111111111111;
20'b01000110000110011101: color_data = 12'b111111111111;
20'b01000110000110011110: color_data = 12'b111111111111;
20'b01000110000110011111: color_data = 12'b111111111111;
20'b01000110000110100000: color_data = 12'b111111111111;
20'b01000110000110100001: color_data = 12'b111111111111;
20'b01000110000110100010: color_data = 12'b111111111111;
20'b01000110000110100011: color_data = 12'b111111111111;
20'b01000110000110100100: color_data = 12'b111111111111;
20'b01000110000110100101: color_data = 12'b111111111111;
20'b01000110000110100110: color_data = 12'b111111111111;
20'b01000110000110100111: color_data = 12'b111111111111;
20'b01000110000110101000: color_data = 12'b111111111111;
20'b01000110000110101001: color_data = 12'b111111111111;
20'b01000110000110101010: color_data = 12'b111111111111;
20'b01000110000110101011: color_data = 12'b111111111111;
20'b01000110000110101100: color_data = 12'b111111111111;
20'b01000110000110101101: color_data = 12'b111111111111;
20'b01000110000110101110: color_data = 12'b111111111111;
20'b01000110000110101111: color_data = 12'b111111111111;
20'b01000110000110110000: color_data = 12'b111111111111;
20'b01000110000110110001: color_data = 12'b111111111111;
20'b01000110000110110010: color_data = 12'b111111111111;
20'b01000110000110110011: color_data = 12'b111111111111;
20'b01000110010011011111: color_data = 12'b111111111111;
20'b01000110010011100000: color_data = 12'b111111111111;
20'b01000110010011100001: color_data = 12'b111111111111;
20'b01000110010011100010: color_data = 12'b111111111111;
20'b01000110010011100011: color_data = 12'b111111111111;
20'b01000110010011100100: color_data = 12'b111111111111;
20'b01000110010011100101: color_data = 12'b111111111111;
20'b01000110010011100110: color_data = 12'b111111111111;
20'b01000110010011100111: color_data = 12'b111111111111;
20'b01000110010011101000: color_data = 12'b111111111111;
20'b01000110010011101001: color_data = 12'b111111111111;
20'b01000110010011110011: color_data = 12'b111111111111;
20'b01000110010011110100: color_data = 12'b111111111111;
20'b01000110010011110101: color_data = 12'b111111111111;
20'b01000110010011110110: color_data = 12'b111111111111;
20'b01000110010011110111: color_data = 12'b111111111111;
20'b01000110010011111000: color_data = 12'b111111111111;
20'b01000110010011111001: color_data = 12'b111111111111;
20'b01000110010011111010: color_data = 12'b111111111111;
20'b01000110010100010101: color_data = 12'b111111111111;
20'b01000110010100010110: color_data = 12'b111111111111;
20'b01000110010100010111: color_data = 12'b111111111111;
20'b01000110010100011000: color_data = 12'b111111111111;
20'b01000110010100011001: color_data = 12'b111111111111;
20'b01000110010100011010: color_data = 12'b111111111111;
20'b01000110010100110100: color_data = 12'b111111111111;
20'b01000110010100110101: color_data = 12'b111111111111;
20'b01000110010100110110: color_data = 12'b111111111111;
20'b01000110010100110111: color_data = 12'b111111111111;
20'b01000110010100111000: color_data = 12'b111111111111;
20'b01000110010100111001: color_data = 12'b111111111111;
20'b01000110010100111010: color_data = 12'b111111111111;
20'b01000110010101001000: color_data = 12'b111111111111;
20'b01000110010101001001: color_data = 12'b111111111111;
20'b01000110010101001010: color_data = 12'b111111111111;
20'b01000110010101001011: color_data = 12'b111111111111;
20'b01000110010101001100: color_data = 12'b111111111111;
20'b01000110010101001101: color_data = 12'b111111111111;
20'b01000110010101010100: color_data = 12'b111111111111;
20'b01000110010101010101: color_data = 12'b111111111111;
20'b01000110010101010110: color_data = 12'b111111111111;
20'b01000110010101010111: color_data = 12'b111111111111;
20'b01000110010101011000: color_data = 12'b111111111111;
20'b01000110010101011001: color_data = 12'b111111111111;
20'b01000110010101011010: color_data = 12'b111111111111;
20'b01000110010101110100: color_data = 12'b111111111111;
20'b01000110010101110101: color_data = 12'b111111111111;
20'b01000110010101110110: color_data = 12'b111111111111;
20'b01000110010101110111: color_data = 12'b111111111111;
20'b01000110010101111000: color_data = 12'b111111111111;
20'b01000110010101111001: color_data = 12'b111111111111;
20'b01000110010110101101: color_data = 12'b111111111111;
20'b01000110010110101110: color_data = 12'b111111111111;
20'b01000110010110101111: color_data = 12'b111111111111;
20'b01000110010110110000: color_data = 12'b111111111111;
20'b01000110010110110001: color_data = 12'b111111111111;
20'b01000110010110110010: color_data = 12'b111111111111;
20'b01000110010110110011: color_data = 12'b111111111111;
20'b01000110100011011111: color_data = 12'b111111111111;
20'b01000110100011100000: color_data = 12'b111111111111;
20'b01000110100011100001: color_data = 12'b111111111111;
20'b01000110100011100010: color_data = 12'b111111111111;
20'b01000110100011100011: color_data = 12'b111111111111;
20'b01000110100011100100: color_data = 12'b111111111111;
20'b01000110100011100101: color_data = 12'b111111111111;
20'b01000110100011100110: color_data = 12'b111111111111;
20'b01000110100011100111: color_data = 12'b111111111111;
20'b01000110100011101000: color_data = 12'b111111111111;
20'b01000110100011101001: color_data = 12'b111111111111;
20'b01000110100011110011: color_data = 12'b111111111111;
20'b01000110100011110100: color_data = 12'b111111111111;
20'b01000110100011110101: color_data = 12'b111111111111;
20'b01000110100011110110: color_data = 12'b111111111111;
20'b01000110100011110111: color_data = 12'b111111111111;
20'b01000110100011111000: color_data = 12'b111111111111;
20'b01000110100011111001: color_data = 12'b111111111111;
20'b01000110100011111010: color_data = 12'b111111111111;
20'b01000110100100010101: color_data = 12'b111111111111;
20'b01000110100100010110: color_data = 12'b111111111111;
20'b01000110100100010111: color_data = 12'b111111111111;
20'b01000110100100011000: color_data = 12'b111111111111;
20'b01000110100100011001: color_data = 12'b111111111111;
20'b01000110100100011010: color_data = 12'b111111111111;
20'b01000110100100110100: color_data = 12'b111111111111;
20'b01000110100100110101: color_data = 12'b111111111111;
20'b01000110100100110110: color_data = 12'b111111111111;
20'b01000110100100110111: color_data = 12'b111111111111;
20'b01000110100100111000: color_data = 12'b111111111111;
20'b01000110100100111001: color_data = 12'b111111111111;
20'b01000110100100111010: color_data = 12'b111111111111;
20'b01000110100101001000: color_data = 12'b111111111111;
20'b01000110100101001001: color_data = 12'b111111111111;
20'b01000110100101001010: color_data = 12'b111111111111;
20'b01000110100101001011: color_data = 12'b111111111111;
20'b01000110100101001100: color_data = 12'b111111111111;
20'b01000110100101001101: color_data = 12'b111111111111;
20'b01000110100101010100: color_data = 12'b111111111111;
20'b01000110100101010101: color_data = 12'b111111111111;
20'b01000110100101010110: color_data = 12'b111111111111;
20'b01000110100101010111: color_data = 12'b111111111111;
20'b01000110100101011000: color_data = 12'b111111111111;
20'b01000110100101011001: color_data = 12'b111111111111;
20'b01000110100101011010: color_data = 12'b111111111111;
20'b01000110100101110100: color_data = 12'b111111111111;
20'b01000110100101110101: color_data = 12'b111111111111;
20'b01000110100101110110: color_data = 12'b111111111111;
20'b01000110100101110111: color_data = 12'b111111111111;
20'b01000110100101111000: color_data = 12'b111111111111;
20'b01000110100101111001: color_data = 12'b111111111111;
20'b01000110100110101101: color_data = 12'b111111111111;
20'b01000110100110101110: color_data = 12'b111111111111;
20'b01000110100110101111: color_data = 12'b111111111111;
20'b01000110100110110000: color_data = 12'b111111111111;
20'b01000110100110110001: color_data = 12'b111111111111;
20'b01000110100110110010: color_data = 12'b111111111111;
20'b01000110100110110011: color_data = 12'b111111111111;
20'b01000110110011011111: color_data = 12'b111111111111;
20'b01000110110011100000: color_data = 12'b111111111111;
20'b01000110110011100001: color_data = 12'b111111111111;
20'b01000110110011100010: color_data = 12'b111111111111;
20'b01000110110011100011: color_data = 12'b111111111111;
20'b01000110110011100100: color_data = 12'b111111111111;
20'b01000110110011100101: color_data = 12'b111111111111;
20'b01000110110011100110: color_data = 12'b111111111111;
20'b01000110110011100111: color_data = 12'b111111111111;
20'b01000110110011101000: color_data = 12'b111111111111;
20'b01000110110011101001: color_data = 12'b111111111111;
20'b01000110110011110011: color_data = 12'b111111111111;
20'b01000110110011110100: color_data = 12'b111111111111;
20'b01000110110011110101: color_data = 12'b111111111111;
20'b01000110110011110110: color_data = 12'b111111111111;
20'b01000110110011110111: color_data = 12'b111111111111;
20'b01000110110011111000: color_data = 12'b111111111111;
20'b01000110110011111001: color_data = 12'b111111111111;
20'b01000110110011111010: color_data = 12'b111111111111;
20'b01000110110100010101: color_data = 12'b111111111111;
20'b01000110110100010110: color_data = 12'b111111111111;
20'b01000110110100010111: color_data = 12'b111111111111;
20'b01000110110100011000: color_data = 12'b111111111111;
20'b01000110110100011001: color_data = 12'b111111111111;
20'b01000110110100011010: color_data = 12'b111111111111;
20'b01000110110100110100: color_data = 12'b111111111111;
20'b01000110110100110101: color_data = 12'b111111111111;
20'b01000110110100110110: color_data = 12'b111111111111;
20'b01000110110100110111: color_data = 12'b111111111111;
20'b01000110110100111000: color_data = 12'b111111111111;
20'b01000110110100111001: color_data = 12'b111111111111;
20'b01000110110100111010: color_data = 12'b111111111111;
20'b01000110110101001000: color_data = 12'b111111111111;
20'b01000110110101001001: color_data = 12'b111111111111;
20'b01000110110101001010: color_data = 12'b111111111111;
20'b01000110110101001011: color_data = 12'b111111111111;
20'b01000110110101001100: color_data = 12'b111111111111;
20'b01000110110101001101: color_data = 12'b111111111111;
20'b01000110110101010100: color_data = 12'b111111111111;
20'b01000110110101010101: color_data = 12'b111111111111;
20'b01000110110101010110: color_data = 12'b111111111111;
20'b01000110110101010111: color_data = 12'b111111111111;
20'b01000110110101011000: color_data = 12'b111111111111;
20'b01000110110101011001: color_data = 12'b111111111111;
20'b01000110110101011010: color_data = 12'b111111111111;
20'b01000110110101110100: color_data = 12'b111111111111;
20'b01000110110101110101: color_data = 12'b111111111111;
20'b01000110110101110110: color_data = 12'b111111111111;
20'b01000110110101110111: color_data = 12'b111111111111;
20'b01000110110101111000: color_data = 12'b111111111111;
20'b01000110110101111001: color_data = 12'b111111111111;
20'b01000110110110101101: color_data = 12'b111111111111;
20'b01000110110110101110: color_data = 12'b111111111111;
20'b01000110110110101111: color_data = 12'b111111111111;
20'b01000110110110110000: color_data = 12'b111111111111;
20'b01000110110110110001: color_data = 12'b111111111111;
20'b01000110110110110010: color_data = 12'b111111111111;
20'b01000110110110110011: color_data = 12'b111111111111;
20'b01000111000011110011: color_data = 12'b111111111111;
20'b01000111000011110100: color_data = 12'b111111111111;
20'b01000111000011110101: color_data = 12'b111111111111;
20'b01000111000011110110: color_data = 12'b111111111111;
20'b01000111000011110111: color_data = 12'b111111111111;
20'b01000111000011111000: color_data = 12'b111111111111;
20'b01000111000011111001: color_data = 12'b111111111111;
20'b01000111000011111010: color_data = 12'b111111111111;
20'b01000111000100010101: color_data = 12'b111111111111;
20'b01000111000100010110: color_data = 12'b111111111111;
20'b01000111000100010111: color_data = 12'b111111111111;
20'b01000111000100011000: color_data = 12'b111111111111;
20'b01000111000100011001: color_data = 12'b111111111111;
20'b01000111000100011010: color_data = 12'b111111111111;
20'b01000111000100110100: color_data = 12'b111111111111;
20'b01000111000100110101: color_data = 12'b111111111111;
20'b01000111000100110110: color_data = 12'b111111111111;
20'b01000111000100110111: color_data = 12'b111111111111;
20'b01000111000100111000: color_data = 12'b111111111111;
20'b01000111000100111001: color_data = 12'b111111111111;
20'b01000111000100111010: color_data = 12'b111111111111;
20'b01000111000101001000: color_data = 12'b111111111111;
20'b01000111000101001001: color_data = 12'b111111111111;
20'b01000111000101001010: color_data = 12'b111111111111;
20'b01000111000101001011: color_data = 12'b111111111111;
20'b01000111000101001100: color_data = 12'b111111111111;
20'b01000111000101001101: color_data = 12'b111111111111;
20'b01000111000101010100: color_data = 12'b111111111111;
20'b01000111000101010101: color_data = 12'b111111111111;
20'b01000111000101010110: color_data = 12'b111111111111;
20'b01000111000101010111: color_data = 12'b111111111111;
20'b01000111000101011000: color_data = 12'b111111111111;
20'b01000111000101011001: color_data = 12'b111111111111;
20'b01000111000101011010: color_data = 12'b111111111111;
20'b01000111000101110100: color_data = 12'b111111111111;
20'b01000111000101110101: color_data = 12'b111111111111;
20'b01000111000101110110: color_data = 12'b111111111111;
20'b01000111000101110111: color_data = 12'b111111111111;
20'b01000111000101111000: color_data = 12'b111111111111;
20'b01000111000101111001: color_data = 12'b111111111111;
20'b01000111000110101101: color_data = 12'b111111111111;
20'b01000111000110101110: color_data = 12'b111111111111;
20'b01000111000110101111: color_data = 12'b111111111111;
20'b01000111000110110000: color_data = 12'b111111111111;
20'b01000111000110110001: color_data = 12'b111111111111;
20'b01000111000110110010: color_data = 12'b111111111111;
20'b01000111000110110011: color_data = 12'b111111111111;
20'b01000111010011110011: color_data = 12'b111111111111;
20'b01000111010011110100: color_data = 12'b111111111111;
20'b01000111010011110101: color_data = 12'b111111111111;
20'b01000111010011110110: color_data = 12'b111111111111;
20'b01000111010011110111: color_data = 12'b111111111111;
20'b01000111010011111000: color_data = 12'b111111111111;
20'b01000111010011111001: color_data = 12'b111111111111;
20'b01000111010011111010: color_data = 12'b111111111111;
20'b01000111010100010101: color_data = 12'b111111111111;
20'b01000111010100010110: color_data = 12'b111111111111;
20'b01000111010100010111: color_data = 12'b111111111111;
20'b01000111010100011000: color_data = 12'b111111111111;
20'b01000111010100011001: color_data = 12'b111111111111;
20'b01000111010100011010: color_data = 12'b111111111111;
20'b01000111010100110100: color_data = 12'b111111111111;
20'b01000111010100110101: color_data = 12'b111111111111;
20'b01000111010100110110: color_data = 12'b111111111111;
20'b01000111010100110111: color_data = 12'b111111111111;
20'b01000111010100111000: color_data = 12'b111111111111;
20'b01000111010100111001: color_data = 12'b111111111111;
20'b01000111010100111010: color_data = 12'b111111111111;
20'b01000111010101001000: color_data = 12'b111111111111;
20'b01000111010101001001: color_data = 12'b111111111111;
20'b01000111010101001010: color_data = 12'b111111111111;
20'b01000111010101001011: color_data = 12'b111111111111;
20'b01000111010101001100: color_data = 12'b111111111111;
20'b01000111010101001101: color_data = 12'b111111111111;
20'b01000111010101010100: color_data = 12'b111111111111;
20'b01000111010101010101: color_data = 12'b111111111111;
20'b01000111010101010110: color_data = 12'b111111111111;
20'b01000111010101010111: color_data = 12'b111111111111;
20'b01000111010101011000: color_data = 12'b111111111111;
20'b01000111010101011001: color_data = 12'b111111111111;
20'b01000111010101011010: color_data = 12'b111111111111;
20'b01000111010101110100: color_data = 12'b111111111111;
20'b01000111010101110101: color_data = 12'b111111111111;
20'b01000111010101110110: color_data = 12'b111111111111;
20'b01000111010101110111: color_data = 12'b111111111111;
20'b01000111010101111000: color_data = 12'b111111111111;
20'b01000111010101111001: color_data = 12'b111111111111;
20'b01000111010110101101: color_data = 12'b111111111111;
20'b01000111010110101110: color_data = 12'b111111111111;
20'b01000111010110101111: color_data = 12'b111111111111;
20'b01000111010110110000: color_data = 12'b111111111111;
20'b01000111010110110001: color_data = 12'b111111111111;
20'b01000111010110110010: color_data = 12'b111111111111;
20'b01000111010110110011: color_data = 12'b111111111111;
20'b01000111100011110011: color_data = 12'b111111111111;
20'b01000111100011110100: color_data = 12'b111111111111;
20'b01000111100011110101: color_data = 12'b111111111111;
20'b01000111100011110110: color_data = 12'b111111111111;
20'b01000111100011110111: color_data = 12'b111111111111;
20'b01000111100011111000: color_data = 12'b111111111111;
20'b01000111100011111001: color_data = 12'b111111111111;
20'b01000111100011111010: color_data = 12'b111111111111;
20'b01000111100100010101: color_data = 12'b111111111111;
20'b01000111100100010110: color_data = 12'b111111111111;
20'b01000111100100010111: color_data = 12'b111111111111;
20'b01000111100100011000: color_data = 12'b111111111111;
20'b01000111100100011001: color_data = 12'b111111111111;
20'b01000111100100011010: color_data = 12'b111111111111;
20'b01000111100100110100: color_data = 12'b111111111111;
20'b01000111100100110101: color_data = 12'b111111111111;
20'b01000111100100110110: color_data = 12'b111111111111;
20'b01000111100100110111: color_data = 12'b111111111111;
20'b01000111100100111000: color_data = 12'b111111111111;
20'b01000111100100111001: color_data = 12'b111111111111;
20'b01000111100100111010: color_data = 12'b111111111111;
20'b01000111100101001000: color_data = 12'b111111111111;
20'b01000111100101001001: color_data = 12'b111111111111;
20'b01000111100101001010: color_data = 12'b111111111111;
20'b01000111100101001011: color_data = 12'b111111111111;
20'b01000111100101001100: color_data = 12'b111111111111;
20'b01000111100101001101: color_data = 12'b111111111111;
20'b01000111100101010100: color_data = 12'b111111111111;
20'b01000111100101010101: color_data = 12'b111111111111;
20'b01000111100101010110: color_data = 12'b111111111111;
20'b01000111100101010111: color_data = 12'b111111111111;
20'b01000111100101011000: color_data = 12'b111111111111;
20'b01000111100101011001: color_data = 12'b111111111111;
20'b01000111100101011010: color_data = 12'b111111111111;
20'b01000111100101110100: color_data = 12'b111111111111;
20'b01000111100101110101: color_data = 12'b111111111111;
20'b01000111100101110110: color_data = 12'b111111111111;
20'b01000111100101110111: color_data = 12'b111111111111;
20'b01000111100101111000: color_data = 12'b111111111111;
20'b01000111100101111001: color_data = 12'b111111111111;
20'b01000111100110101101: color_data = 12'b111111111111;
20'b01000111100110101110: color_data = 12'b111111111111;
20'b01000111100110101111: color_data = 12'b111111111111;
20'b01000111100110110000: color_data = 12'b111111111111;
20'b01000111100110110001: color_data = 12'b111111111111;
20'b01000111100110110010: color_data = 12'b111111111111;
20'b01000111100110110011: color_data = 12'b111111111111;
20'b01000111110011110011: color_data = 12'b111111111111;
20'b01000111110011110100: color_data = 12'b111111111111;
20'b01000111110011110101: color_data = 12'b111111111111;
20'b01000111110011110110: color_data = 12'b111111111111;
20'b01000111110011110111: color_data = 12'b111111111111;
20'b01000111110011111000: color_data = 12'b111111111111;
20'b01000111110011111001: color_data = 12'b111111111111;
20'b01000111110011111010: color_data = 12'b111111111111;
20'b01000111110011111011: color_data = 12'b111111111111;
20'b01000111110011111100: color_data = 12'b111111111111;
20'b01000111110011111101: color_data = 12'b111111111111;
20'b01000111110011111110: color_data = 12'b111111111111;
20'b01000111110011111111: color_data = 12'b111111111111;
20'b01000111110100000000: color_data = 12'b111111111111;
20'b01000111110100000001: color_data = 12'b111111111111;
20'b01000111110100000010: color_data = 12'b111111111111;
20'b01000111110100000011: color_data = 12'b111111111111;
20'b01000111110100000100: color_data = 12'b111111111111;
20'b01000111110100000101: color_data = 12'b111111111111;
20'b01000111110100000110: color_data = 12'b111111111111;
20'b01000111110100000111: color_data = 12'b111111111111;
20'b01000111110100001000: color_data = 12'b111111111111;
20'b01000111110100001001: color_data = 12'b111111111111;
20'b01000111110100001010: color_data = 12'b111111111111;
20'b01000111110100001011: color_data = 12'b111111111111;
20'b01000111110100001100: color_data = 12'b111111111111;
20'b01000111110100001101: color_data = 12'b111111111111;
20'b01000111110100010101: color_data = 12'b111111111111;
20'b01000111110100010110: color_data = 12'b111111111111;
20'b01000111110100010111: color_data = 12'b111111111111;
20'b01000111110100011000: color_data = 12'b111111111111;
20'b01000111110100011001: color_data = 12'b111111111111;
20'b01000111110100011010: color_data = 12'b111111111111;
20'b01000111110100011011: color_data = 12'b111111111111;
20'b01000111110100011100: color_data = 12'b111111111111;
20'b01000111110100011101: color_data = 12'b111111111111;
20'b01000111110100011110: color_data = 12'b111111111111;
20'b01000111110100011111: color_data = 12'b111111111111;
20'b01000111110100100000: color_data = 12'b111111111111;
20'b01000111110100100001: color_data = 12'b111111111111;
20'b01000111110100100010: color_data = 12'b111111111111;
20'b01000111110100100011: color_data = 12'b111111111111;
20'b01000111110100100100: color_data = 12'b111111111111;
20'b01000111110100100101: color_data = 12'b111111111111;
20'b01000111110100100110: color_data = 12'b111111111111;
20'b01000111110100100111: color_data = 12'b111111111111;
20'b01000111110100101000: color_data = 12'b111111111111;
20'b01000111110100101001: color_data = 12'b111111111111;
20'b01000111110100101010: color_data = 12'b111111111111;
20'b01000111110100101011: color_data = 12'b111111111111;
20'b01000111110100101100: color_data = 12'b111111111111;
20'b01000111110100101101: color_data = 12'b111111111111;
20'b01000111110100110100: color_data = 12'b111111111111;
20'b01000111110100110101: color_data = 12'b111111111111;
20'b01000111110100110110: color_data = 12'b111111111111;
20'b01000111110100110111: color_data = 12'b111111111111;
20'b01000111110100111000: color_data = 12'b111111111111;
20'b01000111110100111001: color_data = 12'b111111111111;
20'b01000111110100111010: color_data = 12'b111111111111;
20'b01000111110100111011: color_data = 12'b111111111111;
20'b01000111110100111100: color_data = 12'b111111111111;
20'b01000111110100111101: color_data = 12'b111111111111;
20'b01000111110100111110: color_data = 12'b111111111111;
20'b01000111110100111111: color_data = 12'b111111111111;
20'b01000111110101000000: color_data = 12'b111111111111;
20'b01000111110101000001: color_data = 12'b111111111111;
20'b01000111110101000010: color_data = 12'b111111111111;
20'b01000111110101000011: color_data = 12'b111111111111;
20'b01000111110101000100: color_data = 12'b111111111111;
20'b01000111110101000101: color_data = 12'b111111111111;
20'b01000111110101000110: color_data = 12'b111111111111;
20'b01000111110101000111: color_data = 12'b111111111111;
20'b01000111110101010100: color_data = 12'b111111111111;
20'b01000111110101010101: color_data = 12'b111111111111;
20'b01000111110101010110: color_data = 12'b111111111111;
20'b01000111110101010111: color_data = 12'b111111111111;
20'b01000111110101011000: color_data = 12'b111111111111;
20'b01000111110101011001: color_data = 12'b111111111111;
20'b01000111110101011010: color_data = 12'b111111111111;
20'b01000111110101011011: color_data = 12'b111111111111;
20'b01000111110101011100: color_data = 12'b111111111111;
20'b01000111110101011101: color_data = 12'b111111111111;
20'b01000111110101011110: color_data = 12'b111111111111;
20'b01000111110101011111: color_data = 12'b111111111111;
20'b01000111110101100000: color_data = 12'b111111111111;
20'b01000111110101100001: color_data = 12'b111111111111;
20'b01000111110101100010: color_data = 12'b111111111111;
20'b01000111110101100011: color_data = 12'b111111111111;
20'b01000111110101100100: color_data = 12'b111111111111;
20'b01000111110101100101: color_data = 12'b111111111111;
20'b01000111110101100110: color_data = 12'b111111111111;
20'b01000111110101100111: color_data = 12'b111111111111;
20'b01000111110101101000: color_data = 12'b111111111111;
20'b01000111110101101001: color_data = 12'b111111111111;
20'b01000111110101101010: color_data = 12'b111111111111;
20'b01000111110101101011: color_data = 12'b111111111111;
20'b01000111110101101100: color_data = 12'b111111111111;
20'b01000111110101101101: color_data = 12'b111111111111;
20'b01000111110101110100: color_data = 12'b111111111111;
20'b01000111110101110101: color_data = 12'b111111111111;
20'b01000111110101110110: color_data = 12'b111111111111;
20'b01000111110101110111: color_data = 12'b111111111111;
20'b01000111110101111000: color_data = 12'b111111111111;
20'b01000111110101111001: color_data = 12'b111111111111;
20'b01000111110101111010: color_data = 12'b111111111111;
20'b01000111110101111011: color_data = 12'b111111111111;
20'b01000111110101111100: color_data = 12'b111111111111;
20'b01000111110101111101: color_data = 12'b111111111111;
20'b01000111110101111110: color_data = 12'b111111111111;
20'b01000111110101111111: color_data = 12'b111111111111;
20'b01000111110110000000: color_data = 12'b111111111111;
20'b01000111110110000001: color_data = 12'b111111111111;
20'b01000111110110000010: color_data = 12'b111111111111;
20'b01000111110110000011: color_data = 12'b111111111111;
20'b01000111110110000100: color_data = 12'b111111111111;
20'b01000111110110000101: color_data = 12'b111111111111;
20'b01000111110110000110: color_data = 12'b111111111111;
20'b01000111110110000111: color_data = 12'b111111111111;
20'b01000111110110001000: color_data = 12'b111111111111;
20'b01000111110110001001: color_data = 12'b111111111111;
20'b01000111110110001010: color_data = 12'b111111111111;
20'b01000111110110001011: color_data = 12'b111111111111;
20'b01000111110110001100: color_data = 12'b111111111111;
20'b01000111110110001101: color_data = 12'b111111111111;
20'b01000111110110011010: color_data = 12'b111111111111;
20'b01000111110110011011: color_data = 12'b111111111111;
20'b01000111110110011100: color_data = 12'b111111111111;
20'b01000111110110011101: color_data = 12'b111111111111;
20'b01000111110110011110: color_data = 12'b111111111111;
20'b01000111110110011111: color_data = 12'b111111111111;
20'b01000111110110100000: color_data = 12'b111111111111;
20'b01000111110110100001: color_data = 12'b111111111111;
20'b01000111110110100010: color_data = 12'b111111111111;
20'b01000111110110100011: color_data = 12'b111111111111;
20'b01000111110110100100: color_data = 12'b111111111111;
20'b01000111110110100101: color_data = 12'b111111111111;
20'b01000111110110100110: color_data = 12'b111111111111;
20'b01000111110110100111: color_data = 12'b111111111111;
20'b01000111110110101000: color_data = 12'b111111111111;
20'b01000111110110101001: color_data = 12'b111111111111;
20'b01000111110110101010: color_data = 12'b111111111111;
20'b01000111110110101011: color_data = 12'b111111111111;
20'b01000111110110101100: color_data = 12'b111111111111;
20'b01000111110110101101: color_data = 12'b111111111111;
20'b01000111110110101110: color_data = 12'b111111111111;
20'b01000111110110101111: color_data = 12'b111111111111;
20'b01000111110110110000: color_data = 12'b111111111111;
20'b01000111110110110001: color_data = 12'b111111111111;
20'b01000111110110110010: color_data = 12'b111111111111;
20'b01000111110110110011: color_data = 12'b111111111111;
20'b01001000000011110011: color_data = 12'b111111111111;
20'b01001000000011110100: color_data = 12'b111111111111;
20'b01001000000011110101: color_data = 12'b111111111111;
20'b01001000000011110110: color_data = 12'b111111111111;
20'b01001000000011110111: color_data = 12'b111111111111;
20'b01001000000011111000: color_data = 12'b111111111111;
20'b01001000000011111001: color_data = 12'b111111111111;
20'b01001000000011111010: color_data = 12'b111111111111;
20'b01001000000011111011: color_data = 12'b111111111111;
20'b01001000000011111100: color_data = 12'b111111111111;
20'b01001000000011111101: color_data = 12'b111111111111;
20'b01001000000011111110: color_data = 12'b111111111111;
20'b01001000000011111111: color_data = 12'b111111111111;
20'b01001000000100000000: color_data = 12'b111111111111;
20'b01001000000100000001: color_data = 12'b111111111111;
20'b01001000000100000010: color_data = 12'b111111111111;
20'b01001000000100000011: color_data = 12'b111111111111;
20'b01001000000100000100: color_data = 12'b111111111111;
20'b01001000000100000101: color_data = 12'b111111111111;
20'b01001000000100000110: color_data = 12'b111111111111;
20'b01001000000100000111: color_data = 12'b111111111111;
20'b01001000000100001000: color_data = 12'b111111111111;
20'b01001000000100001001: color_data = 12'b111111111111;
20'b01001000000100001010: color_data = 12'b111111111111;
20'b01001000000100001011: color_data = 12'b111111111111;
20'b01001000000100001100: color_data = 12'b111111111111;
20'b01001000000100001101: color_data = 12'b111111111111;
20'b01001000000100010101: color_data = 12'b111111111111;
20'b01001000000100010110: color_data = 12'b111111111111;
20'b01001000000100010111: color_data = 12'b111111111111;
20'b01001000000100011000: color_data = 12'b111111111111;
20'b01001000000100011001: color_data = 12'b111111111111;
20'b01001000000100011010: color_data = 12'b111111111111;
20'b01001000000100011011: color_data = 12'b111111111111;
20'b01001000000100011100: color_data = 12'b111111111111;
20'b01001000000100011101: color_data = 12'b111111111111;
20'b01001000000100011110: color_data = 12'b111111111111;
20'b01001000000100011111: color_data = 12'b111111111111;
20'b01001000000100100000: color_data = 12'b111111111111;
20'b01001000000100100001: color_data = 12'b111111111111;
20'b01001000000100100010: color_data = 12'b111111111111;
20'b01001000000100100011: color_data = 12'b111111111111;
20'b01001000000100100100: color_data = 12'b111111111111;
20'b01001000000100100101: color_data = 12'b111111111111;
20'b01001000000100100110: color_data = 12'b111111111111;
20'b01001000000100100111: color_data = 12'b111111111111;
20'b01001000000100101000: color_data = 12'b111111111111;
20'b01001000000100101001: color_data = 12'b111111111111;
20'b01001000000100101010: color_data = 12'b111111111111;
20'b01001000000100101011: color_data = 12'b111111111111;
20'b01001000000100101100: color_data = 12'b111111111111;
20'b01001000000100101101: color_data = 12'b111111111111;
20'b01001000000100110100: color_data = 12'b111111111111;
20'b01001000000100110101: color_data = 12'b111111111111;
20'b01001000000100110110: color_data = 12'b111111111111;
20'b01001000000100110111: color_data = 12'b111111111111;
20'b01001000000100111000: color_data = 12'b111111111111;
20'b01001000000100111001: color_data = 12'b111111111111;
20'b01001000000100111010: color_data = 12'b111111111111;
20'b01001000000100111011: color_data = 12'b111111111111;
20'b01001000000100111100: color_data = 12'b111111111111;
20'b01001000000100111101: color_data = 12'b111111111111;
20'b01001000000100111110: color_data = 12'b111111111111;
20'b01001000000100111111: color_data = 12'b111111111111;
20'b01001000000101000000: color_data = 12'b111111111111;
20'b01001000000101000001: color_data = 12'b111111111111;
20'b01001000000101000010: color_data = 12'b111111111111;
20'b01001000000101000011: color_data = 12'b111111111111;
20'b01001000000101000100: color_data = 12'b111111111111;
20'b01001000000101000101: color_data = 12'b111111111111;
20'b01001000000101000110: color_data = 12'b111111111111;
20'b01001000000101000111: color_data = 12'b111111111111;
20'b01001000000101010100: color_data = 12'b111111111111;
20'b01001000000101010101: color_data = 12'b111111111111;
20'b01001000000101010110: color_data = 12'b111111111111;
20'b01001000000101010111: color_data = 12'b111111111111;
20'b01001000000101011000: color_data = 12'b111111111111;
20'b01001000000101011001: color_data = 12'b111111111111;
20'b01001000000101011010: color_data = 12'b111111111111;
20'b01001000000101011011: color_data = 12'b111111111111;
20'b01001000000101011100: color_data = 12'b111111111111;
20'b01001000000101011101: color_data = 12'b111111111111;
20'b01001000000101011110: color_data = 12'b111111111111;
20'b01001000000101011111: color_data = 12'b111111111111;
20'b01001000000101100000: color_data = 12'b111111111111;
20'b01001000000101100001: color_data = 12'b111111111111;
20'b01001000000101100010: color_data = 12'b111111111111;
20'b01001000000101100011: color_data = 12'b111111111111;
20'b01001000000101100100: color_data = 12'b111111111111;
20'b01001000000101100101: color_data = 12'b111111111111;
20'b01001000000101100110: color_data = 12'b111111111111;
20'b01001000000101100111: color_data = 12'b111111111111;
20'b01001000000101101000: color_data = 12'b111111111111;
20'b01001000000101101001: color_data = 12'b111111111111;
20'b01001000000101101010: color_data = 12'b111111111111;
20'b01001000000101101011: color_data = 12'b111111111111;
20'b01001000000101101100: color_data = 12'b111111111111;
20'b01001000000101101101: color_data = 12'b111111111111;
20'b01001000000101110100: color_data = 12'b111111111111;
20'b01001000000101110101: color_data = 12'b111111111111;
20'b01001000000101110110: color_data = 12'b111111111111;
20'b01001000000101110111: color_data = 12'b111111111111;
20'b01001000000101111000: color_data = 12'b111111111111;
20'b01001000000101111001: color_data = 12'b111111111111;
20'b01001000000101111010: color_data = 12'b111111111111;
20'b01001000000101111011: color_data = 12'b111111111111;
20'b01001000000101111100: color_data = 12'b111111111111;
20'b01001000000101111101: color_data = 12'b111111111111;
20'b01001000000101111110: color_data = 12'b111111111111;
20'b01001000000101111111: color_data = 12'b111111111111;
20'b01001000000110000000: color_data = 12'b111111111111;
20'b01001000000110000001: color_data = 12'b111111111111;
20'b01001000000110000010: color_data = 12'b111111111111;
20'b01001000000110000011: color_data = 12'b111111111111;
20'b01001000000110000100: color_data = 12'b111111111111;
20'b01001000000110000101: color_data = 12'b111111111111;
20'b01001000000110000110: color_data = 12'b111111111111;
20'b01001000000110000111: color_data = 12'b111111111111;
20'b01001000000110001000: color_data = 12'b111111111111;
20'b01001000000110001001: color_data = 12'b111111111111;
20'b01001000000110001010: color_data = 12'b111111111111;
20'b01001000000110001011: color_data = 12'b111111111111;
20'b01001000000110001100: color_data = 12'b111111111111;
20'b01001000000110001101: color_data = 12'b111111111111;
20'b01001000000110011010: color_data = 12'b111111111111;
20'b01001000000110011011: color_data = 12'b111111111111;
20'b01001000000110011100: color_data = 12'b111111111111;
20'b01001000000110011101: color_data = 12'b111111111111;
20'b01001000000110011110: color_data = 12'b111111111111;
20'b01001000000110011111: color_data = 12'b111111111111;
20'b01001000000110100000: color_data = 12'b111111111111;
20'b01001000000110100001: color_data = 12'b111111111111;
20'b01001000000110100010: color_data = 12'b111111111111;
20'b01001000000110100011: color_data = 12'b111111111111;
20'b01001000000110100100: color_data = 12'b111111111111;
20'b01001000000110100101: color_data = 12'b111111111111;
20'b01001000000110100110: color_data = 12'b111111111111;
20'b01001000000110100111: color_data = 12'b111111111111;
20'b01001000000110101000: color_data = 12'b111111111111;
20'b01001000000110101001: color_data = 12'b111111111111;
20'b01001000000110101010: color_data = 12'b111111111111;
20'b01001000000110101011: color_data = 12'b111111111111;
20'b01001000000110101100: color_data = 12'b111111111111;
20'b01001000000110101101: color_data = 12'b111111111111;
20'b01001000000110101110: color_data = 12'b111111111111;
20'b01001000000110101111: color_data = 12'b111111111111;
20'b01001000000110110000: color_data = 12'b111111111111;
20'b01001000000110110001: color_data = 12'b111111111111;
20'b01001000000110110010: color_data = 12'b111111111111;
20'b01001000000110110011: color_data = 12'b111111111111;
20'b01001000010011110011: color_data = 12'b111111111111;
20'b01001000010011110100: color_data = 12'b111111111111;
20'b01001000010011110101: color_data = 12'b111111111111;
20'b01001000010011110110: color_data = 12'b111111111111;
20'b01001000010011110111: color_data = 12'b111111111111;
20'b01001000010011111000: color_data = 12'b111111111111;
20'b01001000010011111001: color_data = 12'b111111111111;
20'b01001000010011111010: color_data = 12'b111111111111;
20'b01001000010011111011: color_data = 12'b111111111111;
20'b01001000010011111100: color_data = 12'b111111111111;
20'b01001000010011111101: color_data = 12'b111111111111;
20'b01001000010011111110: color_data = 12'b111111111111;
20'b01001000010011111111: color_data = 12'b111111111111;
20'b01001000010100000000: color_data = 12'b111111111111;
20'b01001000010100000001: color_data = 12'b111111111111;
20'b01001000010100000010: color_data = 12'b111111111111;
20'b01001000010100000011: color_data = 12'b111111111111;
20'b01001000010100000100: color_data = 12'b111111111111;
20'b01001000010100000101: color_data = 12'b111111111111;
20'b01001000010100000110: color_data = 12'b111111111111;
20'b01001000010100000111: color_data = 12'b111111111111;
20'b01001000010100001000: color_data = 12'b111111111111;
20'b01001000010100001001: color_data = 12'b111111111111;
20'b01001000010100001010: color_data = 12'b111111111111;
20'b01001000010100001011: color_data = 12'b111111111111;
20'b01001000010100001100: color_data = 12'b111111111111;
20'b01001000010100001101: color_data = 12'b111111111111;
20'b01001000010100010101: color_data = 12'b111111111111;
20'b01001000010100010110: color_data = 12'b111111111111;
20'b01001000010100010111: color_data = 12'b111111111111;
20'b01001000010100011000: color_data = 12'b111111111111;
20'b01001000010100011001: color_data = 12'b111111111111;
20'b01001000010100011010: color_data = 12'b111111111111;
20'b01001000010100011011: color_data = 12'b111111111111;
20'b01001000010100011100: color_data = 12'b111111111111;
20'b01001000010100011101: color_data = 12'b111111111111;
20'b01001000010100011110: color_data = 12'b111111111111;
20'b01001000010100011111: color_data = 12'b111111111111;
20'b01001000010100100000: color_data = 12'b111111111111;
20'b01001000010100100001: color_data = 12'b111111111111;
20'b01001000010100100010: color_data = 12'b111111111111;
20'b01001000010100100011: color_data = 12'b111111111111;
20'b01001000010100100100: color_data = 12'b111111111111;
20'b01001000010100100101: color_data = 12'b111111111111;
20'b01001000010100100110: color_data = 12'b111111111111;
20'b01001000010100100111: color_data = 12'b111111111111;
20'b01001000010100101000: color_data = 12'b111111111111;
20'b01001000010100101001: color_data = 12'b111111111111;
20'b01001000010100101010: color_data = 12'b111111111111;
20'b01001000010100101011: color_data = 12'b111111111111;
20'b01001000010100101100: color_data = 12'b111111111111;
20'b01001000010100101101: color_data = 12'b111111111111;
20'b01001000010100110100: color_data = 12'b111111111111;
20'b01001000010100110101: color_data = 12'b111111111111;
20'b01001000010100110110: color_data = 12'b111111111111;
20'b01001000010100110111: color_data = 12'b111111111111;
20'b01001000010100111000: color_data = 12'b111111111111;
20'b01001000010100111001: color_data = 12'b111111111111;
20'b01001000010100111010: color_data = 12'b111111111111;
20'b01001000010100111011: color_data = 12'b111111111111;
20'b01001000010100111100: color_data = 12'b111111111111;
20'b01001000010100111101: color_data = 12'b111111111111;
20'b01001000010100111110: color_data = 12'b111111111111;
20'b01001000010100111111: color_data = 12'b111111111111;
20'b01001000010101000000: color_data = 12'b111111111111;
20'b01001000010101000001: color_data = 12'b111111111111;
20'b01001000010101000010: color_data = 12'b111111111111;
20'b01001000010101000011: color_data = 12'b111111111111;
20'b01001000010101000100: color_data = 12'b111111111111;
20'b01001000010101000101: color_data = 12'b111111111111;
20'b01001000010101000110: color_data = 12'b111111111111;
20'b01001000010101000111: color_data = 12'b111111111111;
20'b01001000010101010100: color_data = 12'b111111111111;
20'b01001000010101010101: color_data = 12'b111111111111;
20'b01001000010101010110: color_data = 12'b111111111111;
20'b01001000010101010111: color_data = 12'b111111111111;
20'b01001000010101011000: color_data = 12'b111111111111;
20'b01001000010101011001: color_data = 12'b111111111111;
20'b01001000010101011010: color_data = 12'b111111111111;
20'b01001000010101011011: color_data = 12'b111111111111;
20'b01001000010101011100: color_data = 12'b111111111111;
20'b01001000010101011101: color_data = 12'b111111111111;
20'b01001000010101011110: color_data = 12'b111111111111;
20'b01001000010101011111: color_data = 12'b111111111111;
20'b01001000010101100000: color_data = 12'b111111111111;
20'b01001000010101100001: color_data = 12'b111111111111;
20'b01001000010101100010: color_data = 12'b111111111111;
20'b01001000010101100011: color_data = 12'b111111111111;
20'b01001000010101100100: color_data = 12'b111111111111;
20'b01001000010101100101: color_data = 12'b111111111111;
20'b01001000010101100110: color_data = 12'b111111111111;
20'b01001000010101100111: color_data = 12'b111111111111;
20'b01001000010101101000: color_data = 12'b111111111111;
20'b01001000010101101001: color_data = 12'b111111111111;
20'b01001000010101101010: color_data = 12'b111111111111;
20'b01001000010101101011: color_data = 12'b111111111111;
20'b01001000010101101100: color_data = 12'b111111111111;
20'b01001000010101101101: color_data = 12'b111111111111;
20'b01001000010101110100: color_data = 12'b111111111111;
20'b01001000010101110101: color_data = 12'b111111111111;
20'b01001000010101110110: color_data = 12'b111111111111;
20'b01001000010101110111: color_data = 12'b111111111111;
20'b01001000010101111000: color_data = 12'b111111111111;
20'b01001000010101111001: color_data = 12'b111111111111;
20'b01001000010101111010: color_data = 12'b111111111111;
20'b01001000010101111011: color_data = 12'b111111111111;
20'b01001000010101111100: color_data = 12'b111111111111;
20'b01001000010101111101: color_data = 12'b111111111111;
20'b01001000010101111110: color_data = 12'b111111111111;
20'b01001000010101111111: color_data = 12'b111111111111;
20'b01001000010110000000: color_data = 12'b111111111111;
20'b01001000010110000001: color_data = 12'b111111111111;
20'b01001000010110000010: color_data = 12'b111111111111;
20'b01001000010110000011: color_data = 12'b111111111111;
20'b01001000010110000100: color_data = 12'b111111111111;
20'b01001000010110000101: color_data = 12'b111111111111;
20'b01001000010110000110: color_data = 12'b111111111111;
20'b01001000010110000111: color_data = 12'b111111111111;
20'b01001000010110001000: color_data = 12'b111111111111;
20'b01001000010110001001: color_data = 12'b111111111111;
20'b01001000010110001010: color_data = 12'b111111111111;
20'b01001000010110001011: color_data = 12'b111111111111;
20'b01001000010110001100: color_data = 12'b111111111111;
20'b01001000010110001101: color_data = 12'b111111111111;
20'b01001000010110011010: color_data = 12'b111111111111;
20'b01001000010110011011: color_data = 12'b111111111111;
20'b01001000010110011100: color_data = 12'b111111111111;
20'b01001000010110011101: color_data = 12'b111111111111;
20'b01001000010110011110: color_data = 12'b111111111111;
20'b01001000010110011111: color_data = 12'b111111111111;
20'b01001000010110100000: color_data = 12'b111111111111;
20'b01001000010110100001: color_data = 12'b111111111111;
20'b01001000010110100010: color_data = 12'b111111111111;
20'b01001000010110100011: color_data = 12'b111111111111;
20'b01001000010110100100: color_data = 12'b111111111111;
20'b01001000010110100101: color_data = 12'b111111111111;
20'b01001000010110100110: color_data = 12'b111111111111;
20'b01001000010110100111: color_data = 12'b111111111111;
20'b01001000010110101000: color_data = 12'b111111111111;
20'b01001000010110101001: color_data = 12'b111111111111;
20'b01001000010110101010: color_data = 12'b111111111111;
20'b01001000010110101011: color_data = 12'b111111111111;
20'b01001000010110101100: color_data = 12'b111111111111;
20'b01001000010110101101: color_data = 12'b111111111111;
20'b01001000010110101110: color_data = 12'b111111111111;
20'b01001000010110101111: color_data = 12'b111111111111;
20'b01001000010110110000: color_data = 12'b111111111111;
20'b01001000010110110001: color_data = 12'b111111111111;
20'b01001000010110110010: color_data = 12'b111111111111;
20'b01001000010110110011: color_data = 12'b111111111111;
20'b01001000100011110011: color_data = 12'b111111111111;
20'b01001000100011110100: color_data = 12'b111111111111;
20'b01001000100011110101: color_data = 12'b111111111111;
20'b01001000100011110110: color_data = 12'b111111111111;
20'b01001000100011110111: color_data = 12'b111111111111;
20'b01001000100011111000: color_data = 12'b111111111111;
20'b01001000100011111001: color_data = 12'b111111111111;
20'b01001000100011111010: color_data = 12'b111111111111;
20'b01001000100011111011: color_data = 12'b111111111111;
20'b01001000100011111100: color_data = 12'b111111111111;
20'b01001000100011111101: color_data = 12'b111111111111;
20'b01001000100011111110: color_data = 12'b111111111111;
20'b01001000100011111111: color_data = 12'b111111111111;
20'b01001000100100000000: color_data = 12'b111111111111;
20'b01001000100100000001: color_data = 12'b111111111111;
20'b01001000100100000010: color_data = 12'b111111111111;
20'b01001000100100000011: color_data = 12'b111111111111;
20'b01001000100100000100: color_data = 12'b111111111111;
20'b01001000100100000101: color_data = 12'b111111111111;
20'b01001000100100000110: color_data = 12'b111111111111;
20'b01001000100100000111: color_data = 12'b111111111111;
20'b01001000100100001000: color_data = 12'b111111111111;
20'b01001000100100001001: color_data = 12'b111111111111;
20'b01001000100100001010: color_data = 12'b111111111111;
20'b01001000100100001011: color_data = 12'b111111111111;
20'b01001000100100001100: color_data = 12'b111111111111;
20'b01001000100100001101: color_data = 12'b111111111111;
20'b01001000100100010101: color_data = 12'b111111111111;
20'b01001000100100010110: color_data = 12'b111111111111;
20'b01001000100100010111: color_data = 12'b111111111111;
20'b01001000100100011000: color_data = 12'b111111111111;
20'b01001000100100011001: color_data = 12'b111111111111;
20'b01001000100100011010: color_data = 12'b111111111111;
20'b01001000100100011011: color_data = 12'b111111111111;
20'b01001000100100011100: color_data = 12'b111111111111;
20'b01001000100100011101: color_data = 12'b111111111111;
20'b01001000100100011110: color_data = 12'b111111111111;
20'b01001000100100011111: color_data = 12'b111111111111;
20'b01001000100100100000: color_data = 12'b111111111111;
20'b01001000100100100001: color_data = 12'b111111111111;
20'b01001000100100100010: color_data = 12'b111111111111;
20'b01001000100100100011: color_data = 12'b111111111111;
20'b01001000100100100100: color_data = 12'b111111111111;
20'b01001000100100100101: color_data = 12'b111111111111;
20'b01001000100100100110: color_data = 12'b111111111111;
20'b01001000100100100111: color_data = 12'b111111111111;
20'b01001000100100101000: color_data = 12'b111111111111;
20'b01001000100100101001: color_data = 12'b111111111111;
20'b01001000100100101010: color_data = 12'b111111111111;
20'b01001000100100101011: color_data = 12'b111111111111;
20'b01001000100100101100: color_data = 12'b111111111111;
20'b01001000100100101101: color_data = 12'b111111111111;
20'b01001000100100110100: color_data = 12'b111111111111;
20'b01001000100100110101: color_data = 12'b111111111111;
20'b01001000100100110110: color_data = 12'b111111111111;
20'b01001000100100110111: color_data = 12'b111111111111;
20'b01001000100100111000: color_data = 12'b111111111111;
20'b01001000100100111001: color_data = 12'b111111111111;
20'b01001000100100111010: color_data = 12'b111111111111;
20'b01001000100100111011: color_data = 12'b111111111111;
20'b01001000100100111100: color_data = 12'b111111111111;
20'b01001000100100111101: color_data = 12'b111111111111;
20'b01001000100100111110: color_data = 12'b111111111111;
20'b01001000100100111111: color_data = 12'b111111111111;
20'b01001000100101000000: color_data = 12'b111111111111;
20'b01001000100101000001: color_data = 12'b111111111111;
20'b01001000100101000010: color_data = 12'b111111111111;
20'b01001000100101000011: color_data = 12'b111111111111;
20'b01001000100101000100: color_data = 12'b111111111111;
20'b01001000100101000101: color_data = 12'b111111111111;
20'b01001000100101000110: color_data = 12'b111111111111;
20'b01001000100101000111: color_data = 12'b111111111111;
20'b01001000100101010100: color_data = 12'b111111111111;
20'b01001000100101010101: color_data = 12'b111111111111;
20'b01001000100101010110: color_data = 12'b111111111111;
20'b01001000100101010111: color_data = 12'b111111111111;
20'b01001000100101011000: color_data = 12'b111111111111;
20'b01001000100101011001: color_data = 12'b111111111111;
20'b01001000100101011010: color_data = 12'b111111111111;
20'b01001000100101011011: color_data = 12'b111111111111;
20'b01001000100101011100: color_data = 12'b111111111111;
20'b01001000100101011101: color_data = 12'b111111111111;
20'b01001000100101011110: color_data = 12'b111111111111;
20'b01001000100101011111: color_data = 12'b111111111111;
20'b01001000100101100000: color_data = 12'b111111111111;
20'b01001000100101100001: color_data = 12'b111111111111;
20'b01001000100101100010: color_data = 12'b111111111111;
20'b01001000100101100011: color_data = 12'b111111111111;
20'b01001000100101100100: color_data = 12'b111111111111;
20'b01001000100101100101: color_data = 12'b111111111111;
20'b01001000100101100110: color_data = 12'b111111111111;
20'b01001000100101100111: color_data = 12'b111111111111;
20'b01001000100101101000: color_data = 12'b111111111111;
20'b01001000100101101001: color_data = 12'b111111111111;
20'b01001000100101101010: color_data = 12'b111111111111;
20'b01001000100101101011: color_data = 12'b111111111111;
20'b01001000100101101100: color_data = 12'b111111111111;
20'b01001000100101101101: color_data = 12'b111111111111;
20'b01001000100101110100: color_data = 12'b111111111111;
20'b01001000100101110101: color_data = 12'b111111111111;
20'b01001000100101110110: color_data = 12'b111111111111;
20'b01001000100101110111: color_data = 12'b111111111111;
20'b01001000100101111000: color_data = 12'b111111111111;
20'b01001000100101111001: color_data = 12'b111111111111;
20'b01001000100101111010: color_data = 12'b111111111111;
20'b01001000100101111011: color_data = 12'b111111111111;
20'b01001000100101111100: color_data = 12'b111111111111;
20'b01001000100101111101: color_data = 12'b111111111111;
20'b01001000100101111110: color_data = 12'b111111111111;
20'b01001000100101111111: color_data = 12'b111111111111;
20'b01001000100110000000: color_data = 12'b111111111111;
20'b01001000100110000001: color_data = 12'b111111111111;
20'b01001000100110000010: color_data = 12'b111111111111;
20'b01001000100110000011: color_data = 12'b111111111111;
20'b01001000100110000100: color_data = 12'b111111111111;
20'b01001000100110000101: color_data = 12'b111111111111;
20'b01001000100110000110: color_data = 12'b111111111111;
20'b01001000100110000111: color_data = 12'b111111111111;
20'b01001000100110001000: color_data = 12'b111111111111;
20'b01001000100110001001: color_data = 12'b111111111111;
20'b01001000100110001010: color_data = 12'b111111111111;
20'b01001000100110001011: color_data = 12'b111111111111;
20'b01001000100110001100: color_data = 12'b111111111111;
20'b01001000100110001101: color_data = 12'b111111111111;
20'b01001000100110011010: color_data = 12'b111111111111;
20'b01001000100110011011: color_data = 12'b111111111111;
20'b01001000100110011100: color_data = 12'b111111111111;
20'b01001000100110011101: color_data = 12'b111111111111;
20'b01001000100110011110: color_data = 12'b111111111111;
20'b01001000100110011111: color_data = 12'b111111111111;
20'b01001000100110100000: color_data = 12'b111111111111;
20'b01001000100110100001: color_data = 12'b111111111111;
20'b01001000100110100010: color_data = 12'b111111111111;
20'b01001000100110100011: color_data = 12'b111111111111;
20'b01001000100110100100: color_data = 12'b111111111111;
20'b01001000100110100101: color_data = 12'b111111111111;
20'b01001000100110100110: color_data = 12'b111111111111;
20'b01001000100110100111: color_data = 12'b111111111111;
20'b01001000100110101000: color_data = 12'b111111111111;
20'b01001000100110101001: color_data = 12'b111111111111;
20'b01001000100110101010: color_data = 12'b111111111111;
20'b01001000100110101011: color_data = 12'b111111111111;
20'b01001000100110101100: color_data = 12'b111111111111;
20'b01001000100110101101: color_data = 12'b111111111111;
20'b01001000100110101110: color_data = 12'b111111111111;
20'b01001000100110101111: color_data = 12'b111111111111;
20'b01001000100110110000: color_data = 12'b111111111111;
20'b01001000100110110001: color_data = 12'b111111111111;
20'b01001000100110110010: color_data = 12'b111111111111;
20'b01001000100110110011: color_data = 12'b111111111111;
20'b01001000110011110011: color_data = 12'b111111111111;
20'b01001000110011110100: color_data = 12'b111111111111;
20'b01001000110011110101: color_data = 12'b111111111111;
20'b01001000110011110110: color_data = 12'b111111111111;
20'b01001000110011110111: color_data = 12'b111111111111;
20'b01001000110011111000: color_data = 12'b111111111111;
20'b01001000110011111001: color_data = 12'b111111111111;
20'b01001000110011111010: color_data = 12'b111111111111;
20'b01001000110011111011: color_data = 12'b111111111111;
20'b01001000110011111100: color_data = 12'b111111111111;
20'b01001000110011111101: color_data = 12'b111111111111;
20'b01001000110011111110: color_data = 12'b111111111111;
20'b01001000110011111111: color_data = 12'b111111111111;
20'b01001000110100000000: color_data = 12'b111111111111;
20'b01001000110100000001: color_data = 12'b111111111111;
20'b01001000110100000010: color_data = 12'b111111111111;
20'b01001000110100000011: color_data = 12'b111111111111;
20'b01001000110100000100: color_data = 12'b111111111111;
20'b01001000110100000101: color_data = 12'b111111111111;
20'b01001000110100000110: color_data = 12'b111111111111;
20'b01001000110100000111: color_data = 12'b111111111111;
20'b01001000110100001000: color_data = 12'b111111111111;
20'b01001000110100001001: color_data = 12'b111111111111;
20'b01001000110100001010: color_data = 12'b111111111111;
20'b01001000110100001011: color_data = 12'b111111111111;
20'b01001000110100001100: color_data = 12'b111111111111;
20'b01001000110100001101: color_data = 12'b111111111111;
20'b01001000110100010101: color_data = 12'b111111111111;
20'b01001000110100010110: color_data = 12'b111111111111;
20'b01001000110100010111: color_data = 12'b111111111111;
20'b01001000110100011000: color_data = 12'b111111111111;
20'b01001000110100011001: color_data = 12'b111111111111;
20'b01001000110100011010: color_data = 12'b111111111111;
20'b01001000110100011011: color_data = 12'b111111111111;
20'b01001000110100011100: color_data = 12'b111111111111;
20'b01001000110100011101: color_data = 12'b111111111111;
20'b01001000110100011110: color_data = 12'b111111111111;
20'b01001000110100011111: color_data = 12'b111111111111;
20'b01001000110100100000: color_data = 12'b111111111111;
20'b01001000110100100001: color_data = 12'b111111111111;
20'b01001000110100100010: color_data = 12'b111111111111;
20'b01001000110100100011: color_data = 12'b111111111111;
20'b01001000110100100100: color_data = 12'b111111111111;
20'b01001000110100100101: color_data = 12'b111111111111;
20'b01001000110100100110: color_data = 12'b111111111111;
20'b01001000110100100111: color_data = 12'b111111111111;
20'b01001000110100101000: color_data = 12'b111111111111;
20'b01001000110100101001: color_data = 12'b111111111111;
20'b01001000110100101010: color_data = 12'b111111111111;
20'b01001000110100101011: color_data = 12'b111111111111;
20'b01001000110100101100: color_data = 12'b111111111111;
20'b01001000110100101101: color_data = 12'b111111111111;
20'b01001000110100110100: color_data = 12'b111111111111;
20'b01001000110100110101: color_data = 12'b111111111111;
20'b01001000110100110110: color_data = 12'b111111111111;
20'b01001000110100110111: color_data = 12'b111111111111;
20'b01001000110100111000: color_data = 12'b111111111111;
20'b01001000110100111001: color_data = 12'b111111111111;
20'b01001000110100111010: color_data = 12'b111111111111;
20'b01001000110100111011: color_data = 12'b111111111111;
20'b01001000110100111100: color_data = 12'b111111111111;
20'b01001000110100111101: color_data = 12'b111111111111;
20'b01001000110100111110: color_data = 12'b111111111111;
20'b01001000110100111111: color_data = 12'b111111111111;
20'b01001000110101000000: color_data = 12'b111111111111;
20'b01001000110101000001: color_data = 12'b111111111111;
20'b01001000110101000010: color_data = 12'b111111111111;
20'b01001000110101000011: color_data = 12'b111111111111;
20'b01001000110101000100: color_data = 12'b111111111111;
20'b01001000110101000101: color_data = 12'b111111111111;
20'b01001000110101000110: color_data = 12'b111111111111;
20'b01001000110101000111: color_data = 12'b111111111111;
20'b01001000110101010100: color_data = 12'b111111111111;
20'b01001000110101010101: color_data = 12'b111111111111;
20'b01001000110101010110: color_data = 12'b111111111111;
20'b01001000110101010111: color_data = 12'b111111111111;
20'b01001000110101011000: color_data = 12'b111111111111;
20'b01001000110101011001: color_data = 12'b111111111111;
20'b01001000110101011010: color_data = 12'b111111111111;
20'b01001000110101011011: color_data = 12'b111111111111;
20'b01001000110101011100: color_data = 12'b111111111111;
20'b01001000110101011101: color_data = 12'b111111111111;
20'b01001000110101011110: color_data = 12'b111111111111;
20'b01001000110101011111: color_data = 12'b111111111111;
20'b01001000110101100000: color_data = 12'b111111111111;
20'b01001000110101100001: color_data = 12'b111111111111;
20'b01001000110101100010: color_data = 12'b111111111111;
20'b01001000110101100011: color_data = 12'b111111111111;
20'b01001000110101100100: color_data = 12'b111111111111;
20'b01001000110101100101: color_data = 12'b111111111111;
20'b01001000110101100110: color_data = 12'b111111111111;
20'b01001000110101100111: color_data = 12'b111111111111;
20'b01001000110101101000: color_data = 12'b111111111111;
20'b01001000110101101001: color_data = 12'b111111111111;
20'b01001000110101101010: color_data = 12'b111111111111;
20'b01001000110101101011: color_data = 12'b111111111111;
20'b01001000110101101100: color_data = 12'b111111111111;
20'b01001000110101101101: color_data = 12'b111111111111;
20'b01001000110101110100: color_data = 12'b111111111111;
20'b01001000110101110101: color_data = 12'b111111111111;
20'b01001000110101110110: color_data = 12'b111111111111;
20'b01001000110101110111: color_data = 12'b111111111111;
20'b01001000110101111000: color_data = 12'b111111111111;
20'b01001000110101111001: color_data = 12'b111111111111;
20'b01001000110101111010: color_data = 12'b111111111111;
20'b01001000110101111011: color_data = 12'b111111111111;
20'b01001000110101111100: color_data = 12'b111111111111;
20'b01001000110101111101: color_data = 12'b111111111111;
20'b01001000110101111110: color_data = 12'b111111111111;
20'b01001000110101111111: color_data = 12'b111111111111;
20'b01001000110110000000: color_data = 12'b111111111111;
20'b01001000110110000001: color_data = 12'b111111111111;
20'b01001000110110000010: color_data = 12'b111111111111;
20'b01001000110110000011: color_data = 12'b111111111111;
20'b01001000110110000100: color_data = 12'b111111111111;
20'b01001000110110000101: color_data = 12'b111111111111;
20'b01001000110110000110: color_data = 12'b111111111111;
20'b01001000110110000111: color_data = 12'b111111111111;
20'b01001000110110001000: color_data = 12'b111111111111;
20'b01001000110110001001: color_data = 12'b111111111111;
20'b01001000110110001010: color_data = 12'b111111111111;
20'b01001000110110001011: color_data = 12'b111111111111;
20'b01001000110110001100: color_data = 12'b111111111111;
20'b01001000110110001101: color_data = 12'b111111111111;
20'b01001000110110011010: color_data = 12'b111111111111;
20'b01001000110110011011: color_data = 12'b111111111111;
20'b01001000110110011100: color_data = 12'b111111111111;
20'b01001000110110011101: color_data = 12'b111111111111;
20'b01001000110110011110: color_data = 12'b111111111111;
20'b01001000110110011111: color_data = 12'b111111111111;
20'b01001000110110100000: color_data = 12'b111111111111;
20'b01001000110110100001: color_data = 12'b111111111111;
20'b01001000110110100010: color_data = 12'b111111111111;
20'b01001000110110100011: color_data = 12'b111111111111;
20'b01001000110110100100: color_data = 12'b111111111111;
20'b01001000110110100101: color_data = 12'b111111111111;
20'b01001000110110100110: color_data = 12'b111111111111;
20'b01001000110110100111: color_data = 12'b111111111111;
20'b01001000110110101000: color_data = 12'b111111111111;
20'b01001000110110101001: color_data = 12'b111111111111;
20'b01001000110110101010: color_data = 12'b111111111111;
20'b01001000110110101011: color_data = 12'b111111111111;
20'b01001000110110101100: color_data = 12'b111111111111;
20'b01001000110110101101: color_data = 12'b111111111111;
20'b01001000110110101110: color_data = 12'b111111111111;
20'b01001000110110101111: color_data = 12'b111111111111;
20'b01001000110110110000: color_data = 12'b111111111111;
20'b01001000110110110001: color_data = 12'b111111111111;
20'b01001000110110110010: color_data = 12'b111111111111;
20'b01001000110110110011: color_data = 12'b111111111111;
20'b01001001000011110011: color_data = 12'b111111111111;
20'b01001001000011110100: color_data = 12'b111111111111;
20'b01001001000011110101: color_data = 12'b111111111111;
20'b01001001000011110110: color_data = 12'b111111111111;
20'b01001001000011110111: color_data = 12'b111111111111;
20'b01001001000011111000: color_data = 12'b111111111111;
20'b01001001000011111001: color_data = 12'b111111111111;
20'b01001001000011111010: color_data = 12'b111111111111;
20'b01001001000011111011: color_data = 12'b111111111111;
20'b01001001000011111100: color_data = 12'b111111111111;
20'b01001001000011111101: color_data = 12'b111111111111;
20'b01001001000011111110: color_data = 12'b111111111111;
20'b01001001000011111111: color_data = 12'b111111111111;
20'b01001001000100000000: color_data = 12'b111111111111;
20'b01001001000100000001: color_data = 12'b111111111111;
20'b01001001000100000010: color_data = 12'b111111111111;
20'b01001001000100000011: color_data = 12'b111111111111;
20'b01001001000100000100: color_data = 12'b111111111111;
20'b01001001000100000101: color_data = 12'b111111111111;
20'b01001001000100000110: color_data = 12'b111111111111;
20'b01001001000100000111: color_data = 12'b111111111111;
20'b01001001000100001000: color_data = 12'b111111111111;
20'b01001001000100001001: color_data = 12'b111111111111;
20'b01001001000100001010: color_data = 12'b111111111111;
20'b01001001000100001011: color_data = 12'b111111111111;
20'b01001001000100001100: color_data = 12'b111111111111;
20'b01001001000100001101: color_data = 12'b111111111111;
20'b01001001000100010101: color_data = 12'b111111111111;
20'b01001001000100010110: color_data = 12'b111111111111;
20'b01001001000100010111: color_data = 12'b111111111111;
20'b01001001000100011000: color_data = 12'b111111111111;
20'b01001001000100011001: color_data = 12'b111111111111;
20'b01001001000100011010: color_data = 12'b111111111111;
20'b01001001000100011011: color_data = 12'b111111111111;
20'b01001001000100011100: color_data = 12'b111111111111;
20'b01001001000100011101: color_data = 12'b111111111111;
20'b01001001000100011110: color_data = 12'b111111111111;
20'b01001001000100011111: color_data = 12'b111111111111;
20'b01001001000100100000: color_data = 12'b111111111111;
20'b01001001000100100001: color_data = 12'b111111111111;
20'b01001001000100100010: color_data = 12'b111111111111;
20'b01001001000100100011: color_data = 12'b111111111111;
20'b01001001000100100100: color_data = 12'b111111111111;
20'b01001001000100100101: color_data = 12'b111111111111;
20'b01001001000100100110: color_data = 12'b111111111111;
20'b01001001000100100111: color_data = 12'b111111111111;
20'b01001001000100101000: color_data = 12'b111111111111;
20'b01001001000100101001: color_data = 12'b111111111111;
20'b01001001000100101010: color_data = 12'b111111111111;
20'b01001001000100101011: color_data = 12'b111111111111;
20'b01001001000100101100: color_data = 12'b111111111111;
20'b01001001000100101101: color_data = 12'b111111111111;
20'b01001001000100110100: color_data = 12'b111111111111;
20'b01001001000100110101: color_data = 12'b111111111111;
20'b01001001000100110110: color_data = 12'b111111111111;
20'b01001001000100110111: color_data = 12'b111111111111;
20'b01001001000100111000: color_data = 12'b111111111111;
20'b01001001000100111001: color_data = 12'b111111111111;
20'b01001001000100111010: color_data = 12'b111111111111;
20'b01001001000100111011: color_data = 12'b111111111111;
20'b01001001000100111100: color_data = 12'b111111111111;
20'b01001001000100111101: color_data = 12'b111111111111;
20'b01001001000100111110: color_data = 12'b111111111111;
20'b01001001000100111111: color_data = 12'b111111111111;
20'b01001001000101000000: color_data = 12'b111111111111;
20'b01001001000101000001: color_data = 12'b111111111111;
20'b01001001000101000010: color_data = 12'b111111111111;
20'b01001001000101000011: color_data = 12'b111111111111;
20'b01001001000101000100: color_data = 12'b111111111111;
20'b01001001000101000101: color_data = 12'b111111111111;
20'b01001001000101000110: color_data = 12'b111111111111;
20'b01001001000101000111: color_data = 12'b111111111111;
20'b01001001000101010100: color_data = 12'b111111111111;
20'b01001001000101010101: color_data = 12'b111111111111;
20'b01001001000101010110: color_data = 12'b111111111111;
20'b01001001000101010111: color_data = 12'b111111111111;
20'b01001001000101011000: color_data = 12'b111111111111;
20'b01001001000101011001: color_data = 12'b111111111111;
20'b01001001000101011010: color_data = 12'b111111111111;
20'b01001001000101011011: color_data = 12'b111111111111;
20'b01001001000101011100: color_data = 12'b111111111111;
20'b01001001000101011101: color_data = 12'b111111111111;
20'b01001001000101011110: color_data = 12'b111111111111;
20'b01001001000101011111: color_data = 12'b111111111111;
20'b01001001000101100000: color_data = 12'b111111111111;
20'b01001001000101100001: color_data = 12'b111111111111;
20'b01001001000101100010: color_data = 12'b111111111111;
20'b01001001000101100011: color_data = 12'b111111111111;
20'b01001001000101100100: color_data = 12'b111111111111;
20'b01001001000101100101: color_data = 12'b111111111111;
20'b01001001000101100110: color_data = 12'b111111111111;
20'b01001001000101100111: color_data = 12'b111111111111;
20'b01001001000101101000: color_data = 12'b111111111111;
20'b01001001000101101001: color_data = 12'b111111111111;
20'b01001001000101101010: color_data = 12'b111111111111;
20'b01001001000101101011: color_data = 12'b111111111111;
20'b01001001000101101100: color_data = 12'b111111111111;
20'b01001001000101101101: color_data = 12'b111111111111;
20'b01001001000101110100: color_data = 12'b111111111111;
20'b01001001000101110101: color_data = 12'b111111111111;
20'b01001001000101110110: color_data = 12'b111111111111;
20'b01001001000101110111: color_data = 12'b111111111111;
20'b01001001000101111000: color_data = 12'b111111111111;
20'b01001001000101111001: color_data = 12'b111111111111;
20'b01001001000101111010: color_data = 12'b111111111111;
20'b01001001000101111011: color_data = 12'b111111111111;
20'b01001001000101111100: color_data = 12'b111111111111;
20'b01001001000101111101: color_data = 12'b111111111111;
20'b01001001000101111110: color_data = 12'b111111111111;
20'b01001001000101111111: color_data = 12'b111111111111;
20'b01001001000110000000: color_data = 12'b111111111111;
20'b01001001000110000001: color_data = 12'b111111111111;
20'b01001001000110000010: color_data = 12'b111111111111;
20'b01001001000110000011: color_data = 12'b111111111111;
20'b01001001000110000100: color_data = 12'b111111111111;
20'b01001001000110000101: color_data = 12'b111111111111;
20'b01001001000110000110: color_data = 12'b111111111111;
20'b01001001000110000111: color_data = 12'b111111111111;
20'b01001001000110001000: color_data = 12'b111111111111;
20'b01001001000110001001: color_data = 12'b111111111111;
20'b01001001000110001010: color_data = 12'b111111111111;
20'b01001001000110001011: color_data = 12'b111111111111;
20'b01001001000110001100: color_data = 12'b111111111111;
20'b01001001000110001101: color_data = 12'b111111111111;
20'b01001001000110011010: color_data = 12'b111111111111;
20'b01001001000110011011: color_data = 12'b111111111111;
20'b01001001000110011100: color_data = 12'b111111111111;
20'b01001001000110011101: color_data = 12'b111111111111;
20'b01001001000110011110: color_data = 12'b111111111111;
20'b01001001000110011111: color_data = 12'b111111111111;
20'b01001001000110100000: color_data = 12'b111111111111;
20'b01001001000110100001: color_data = 12'b111111111111;
20'b01001001000110100010: color_data = 12'b111111111111;
20'b01001001000110100011: color_data = 12'b111111111111;
20'b01001001000110100100: color_data = 12'b111111111111;
20'b01001001000110100101: color_data = 12'b111111111111;
20'b01001001000110100110: color_data = 12'b111111111111;
20'b01001001000110100111: color_data = 12'b111111111111;
20'b01001001000110101000: color_data = 12'b111111111111;
20'b01001001000110101001: color_data = 12'b111111111111;
20'b01001001000110101010: color_data = 12'b111111111111;
20'b01001001000110101011: color_data = 12'b111111111111;
20'b01001001000110101100: color_data = 12'b111111111111;
20'b01001001000110101101: color_data = 12'b111111111111;
20'b01001001000110101110: color_data = 12'b111111111111;
20'b01001001000110101111: color_data = 12'b111111111111;
20'b01001001000110110000: color_data = 12'b111111111111;
20'b01001001000110110001: color_data = 12'b111111111111;
20'b01001001000110110010: color_data = 12'b111111111111;
20'b01001001000110110011: color_data = 12'b111111111111;
20'b01001001010011110011: color_data = 12'b111111111111;
20'b01001001010011110100: color_data = 12'b111111111111;
20'b01001001010011110101: color_data = 12'b111111111111;
20'b01001001010011110110: color_data = 12'b111111111111;
20'b01001001010011110111: color_data = 12'b111111111111;
20'b01001001010011111000: color_data = 12'b111111111111;
20'b01001001010011111001: color_data = 12'b111111111111;
20'b01001001010011111010: color_data = 12'b111111111111;
20'b01001001010011111011: color_data = 12'b111111111111;
20'b01001001010011111100: color_data = 12'b111111111111;
20'b01001001010011111101: color_data = 12'b111111111111;
20'b01001001010011111110: color_data = 12'b111111111111;
20'b01001001010011111111: color_data = 12'b111111111111;
20'b01001001010100000000: color_data = 12'b111111111111;
20'b01001001010100000001: color_data = 12'b111111111111;
20'b01001001010100000010: color_data = 12'b111111111111;
20'b01001001010100000011: color_data = 12'b111111111111;
20'b01001001010100000100: color_data = 12'b111111111111;
20'b01001001010100000101: color_data = 12'b111111111111;
20'b01001001010100000110: color_data = 12'b111111111111;
20'b01001001010100000111: color_data = 12'b111111111111;
20'b01001001010100001000: color_data = 12'b111111111111;
20'b01001001010100001001: color_data = 12'b111111111111;
20'b01001001010100001010: color_data = 12'b111111111111;
20'b01001001010100001011: color_data = 12'b111111111111;
20'b01001001010100001100: color_data = 12'b111111111111;
20'b01001001010100001101: color_data = 12'b111111111111;
20'b01001001010100010101: color_data = 12'b111111111111;
20'b01001001010100010110: color_data = 12'b111111111111;
20'b01001001010100010111: color_data = 12'b111111111111;
20'b01001001010100011000: color_data = 12'b111111111111;
20'b01001001010100011001: color_data = 12'b111111111111;
20'b01001001010100011010: color_data = 12'b111111111111;
20'b01001001010100011011: color_data = 12'b111111111111;
20'b01001001010100011100: color_data = 12'b111111111111;
20'b01001001010100011101: color_data = 12'b111111111111;
20'b01001001010100011110: color_data = 12'b111111111111;
20'b01001001010100011111: color_data = 12'b111111111111;
20'b01001001010100100000: color_data = 12'b111111111111;
20'b01001001010100100001: color_data = 12'b111111111111;
20'b01001001010100100010: color_data = 12'b111111111111;
20'b01001001010100100011: color_data = 12'b111111111111;
20'b01001001010100100100: color_data = 12'b111111111111;
20'b01001001010100100101: color_data = 12'b111111111111;
20'b01001001010100100110: color_data = 12'b111111111111;
20'b01001001010100100111: color_data = 12'b111111111111;
20'b01001001010100101000: color_data = 12'b111111111111;
20'b01001001010100101001: color_data = 12'b111111111111;
20'b01001001010100101010: color_data = 12'b111111111111;
20'b01001001010100101011: color_data = 12'b111111111111;
20'b01001001010100101100: color_data = 12'b111111111111;
20'b01001001010100101101: color_data = 12'b111111111111;
20'b01001001010100110100: color_data = 12'b111111111111;
20'b01001001010100110101: color_data = 12'b111111111111;
20'b01001001010100110110: color_data = 12'b111111111111;
20'b01001001010100110111: color_data = 12'b111111111111;
20'b01001001010100111000: color_data = 12'b111111111111;
20'b01001001010100111001: color_data = 12'b111111111111;
20'b01001001010100111010: color_data = 12'b111111111111;
20'b01001001010100111011: color_data = 12'b111111111111;
20'b01001001010100111100: color_data = 12'b111111111111;
20'b01001001010100111101: color_data = 12'b111111111111;
20'b01001001010100111110: color_data = 12'b111111111111;
20'b01001001010100111111: color_data = 12'b111111111111;
20'b01001001010101000000: color_data = 12'b111111111111;
20'b01001001010101000001: color_data = 12'b111111111111;
20'b01001001010101000010: color_data = 12'b111111111111;
20'b01001001010101000011: color_data = 12'b111111111111;
20'b01001001010101000100: color_data = 12'b111111111111;
20'b01001001010101000101: color_data = 12'b111111111111;
20'b01001001010101000110: color_data = 12'b111111111111;
20'b01001001010101000111: color_data = 12'b111111111111;
20'b01001001010101010100: color_data = 12'b111111111111;
20'b01001001010101010101: color_data = 12'b111111111111;
20'b01001001010101010110: color_data = 12'b111111111111;
20'b01001001010101010111: color_data = 12'b111111111111;
20'b01001001010101011000: color_data = 12'b111111111111;
20'b01001001010101011001: color_data = 12'b111111111111;
20'b01001001010101011010: color_data = 12'b111111111111;
20'b01001001010101011011: color_data = 12'b111111111111;
20'b01001001010101011100: color_data = 12'b111111111111;
20'b01001001010101011101: color_data = 12'b111111111111;
20'b01001001010101011110: color_data = 12'b111111111111;
20'b01001001010101011111: color_data = 12'b111111111111;
20'b01001001010101100000: color_data = 12'b111111111111;
20'b01001001010101100001: color_data = 12'b111111111111;
20'b01001001010101100010: color_data = 12'b111111111111;
20'b01001001010101100011: color_data = 12'b111111111111;
20'b01001001010101100100: color_data = 12'b111111111111;
20'b01001001010101100101: color_data = 12'b111111111111;
20'b01001001010101100110: color_data = 12'b111111111111;
20'b01001001010101100111: color_data = 12'b111111111111;
20'b01001001010101101000: color_data = 12'b111111111111;
20'b01001001010101101001: color_data = 12'b111111111111;
20'b01001001010101101010: color_data = 12'b111111111111;
20'b01001001010101101011: color_data = 12'b111111111111;
20'b01001001010101101100: color_data = 12'b111111111111;
20'b01001001010101101101: color_data = 12'b111111111111;
20'b01001001010101110100: color_data = 12'b111111111111;
20'b01001001010101110101: color_data = 12'b111111111111;
20'b01001001010101110110: color_data = 12'b111111111111;
20'b01001001010101110111: color_data = 12'b111111111111;
20'b01001001010101111000: color_data = 12'b111111111111;
20'b01001001010101111001: color_data = 12'b111111111111;
20'b01001001010101111010: color_data = 12'b111111111111;
20'b01001001010101111011: color_data = 12'b111111111111;
20'b01001001010101111100: color_data = 12'b111111111111;
20'b01001001010101111101: color_data = 12'b111111111111;
20'b01001001010101111110: color_data = 12'b111111111111;
20'b01001001010101111111: color_data = 12'b111111111111;
20'b01001001010110000000: color_data = 12'b111111111111;
20'b01001001010110000001: color_data = 12'b111111111111;
20'b01001001010110000010: color_data = 12'b111111111111;
20'b01001001010110000011: color_data = 12'b111111111111;
20'b01001001010110000100: color_data = 12'b111111111111;
20'b01001001010110000101: color_data = 12'b111111111111;
20'b01001001010110000110: color_data = 12'b111111111111;
20'b01001001010110000111: color_data = 12'b111111111111;
20'b01001001010110001000: color_data = 12'b111111111111;
20'b01001001010110001001: color_data = 12'b111111111111;
20'b01001001010110001010: color_data = 12'b111111111111;
20'b01001001010110001011: color_data = 12'b111111111111;
20'b01001001010110001100: color_data = 12'b111111111111;
20'b01001001010110001101: color_data = 12'b111111111111;
20'b01001001010110011010: color_data = 12'b111111111111;
20'b01001001010110011011: color_data = 12'b111111111111;
20'b01001001010110011100: color_data = 12'b111111111111;
20'b01001001010110011101: color_data = 12'b111111111111;
20'b01001001010110011110: color_data = 12'b111111111111;
20'b01001001010110011111: color_data = 12'b111111111111;
20'b01001001010110100000: color_data = 12'b111111111111;
20'b01001001010110100001: color_data = 12'b111111111111;
20'b01001001010110100010: color_data = 12'b111111111111;
20'b01001001010110100011: color_data = 12'b111111111111;
20'b01001001010110100100: color_data = 12'b111111111111;
20'b01001001010110100101: color_data = 12'b111111111111;
20'b01001001010110100110: color_data = 12'b111111111111;
20'b01001001010110100111: color_data = 12'b111111111111;
20'b01001001010110101000: color_data = 12'b111111111111;
20'b01001001010110101001: color_data = 12'b111111111111;
20'b01001001010110101010: color_data = 12'b111111111111;
20'b01001001010110101011: color_data = 12'b111111111111;
20'b01001001010110101100: color_data = 12'b111111111111;
20'b01001001010110101101: color_data = 12'b111111111111;
20'b01001001010110101110: color_data = 12'b111111111111;
20'b01001001010110101111: color_data = 12'b111111111111;
20'b01001001010110110000: color_data = 12'b111111111111;
20'b01001001010110110001: color_data = 12'b111111111111;
20'b01001001010110110010: color_data = 12'b111111111111;
20'b01001001010110110011: color_data = 12'b111111111111;
20'b01011001100011111010: color_data = 12'b000011111111;
20'b01011001100011111011: color_data = 12'b000011111111;
20'b01011001100011111100: color_data = 12'b000011111111;
20'b01011001100011111101: color_data = 12'b000011111111;
20'b01011001100011111110: color_data = 12'b000011111111;
20'b01011001100011111111: color_data = 12'b000011111111;
20'b01011001100100000000: color_data = 12'b000011111111;
20'b01011001100100000001: color_data = 12'b000011111111;
20'b01011001100100000010: color_data = 12'b000011111111;
20'b01011001100100000011: color_data = 12'b000011111111;
20'b01011001100100000100: color_data = 12'b000011111111;
20'b01011001100100000101: color_data = 12'b000011111111;
20'b01011001100100000110: color_data = 12'b000011111111;
20'b01011001100100000111: color_data = 12'b000011111111;
20'b01011001100100001000: color_data = 12'b000011111111;
20'b01011001100100001001: color_data = 12'b000011111111;
20'b01011001100100001010: color_data = 12'b000011111111;
20'b01011001100100001011: color_data = 12'b000011111111;
20'b01011001100100001111: color_data = 12'b000011111111;
20'b01011001100100010000: color_data = 12'b000011111111;
20'b01011001100100010001: color_data = 12'b000011111111;
20'b01011001100100010010: color_data = 12'b000011111111;
20'b01011001100100010011: color_data = 12'b000011111111;
20'b01011001100100010100: color_data = 12'b000011111111;
20'b01011001100100010101: color_data = 12'b000011111111;
20'b01011001100100010110: color_data = 12'b000011111111;
20'b01011001100100010111: color_data = 12'b000011111111;
20'b01011001100100011000: color_data = 12'b000011111111;
20'b01011001100100011001: color_data = 12'b000011111111;
20'b01011001100100011010: color_data = 12'b000011111111;
20'b01011001100100011011: color_data = 12'b000011111111;
20'b01011001100100011100: color_data = 12'b000011111111;
20'b01011001100100011101: color_data = 12'b000011111111;
20'b01011001100100011110: color_data = 12'b000011111111;
20'b01011001100100011111: color_data = 12'b000011111111;
20'b01011001100100100000: color_data = 12'b000011111111;
20'b01011001110011111010: color_data = 12'b000011111111;
20'b01011001110011111011: color_data = 12'b000011111111;
20'b01011001110011111100: color_data = 12'b000011111111;
20'b01011001110011111101: color_data = 12'b000011111111;
20'b01011001110011111110: color_data = 12'b000011111111;
20'b01011001110011111111: color_data = 12'b000011111111;
20'b01011001110100000000: color_data = 12'b000011111111;
20'b01011001110100000001: color_data = 12'b000011111111;
20'b01011001110100000010: color_data = 12'b000011111111;
20'b01011001110100000011: color_data = 12'b000011111111;
20'b01011001110100000100: color_data = 12'b000011111111;
20'b01011001110100000101: color_data = 12'b000011111111;
20'b01011001110100000110: color_data = 12'b000011111111;
20'b01011001110100000111: color_data = 12'b000011111111;
20'b01011001110100001000: color_data = 12'b000011111111;
20'b01011001110100001001: color_data = 12'b000011111111;
20'b01011001110100001010: color_data = 12'b000011111111;
20'b01011001110100001011: color_data = 12'b000011111111;
20'b01011001110100001111: color_data = 12'b000011111111;
20'b01011001110100010000: color_data = 12'b000011111111;
20'b01011001110100010001: color_data = 12'b000011111111;
20'b01011001110100010010: color_data = 12'b000011111111;
20'b01011001110100010011: color_data = 12'b000011111111;
20'b01011001110100010100: color_data = 12'b000011111111;
20'b01011001110100010101: color_data = 12'b000011111111;
20'b01011001110100010110: color_data = 12'b000011111111;
20'b01011001110100010111: color_data = 12'b000011111111;
20'b01011001110100011000: color_data = 12'b000011111111;
20'b01011001110100011001: color_data = 12'b000011111111;
20'b01011001110100011010: color_data = 12'b000011111111;
20'b01011001110100011011: color_data = 12'b000011111111;
20'b01011001110100011100: color_data = 12'b000011111111;
20'b01011001110100011101: color_data = 12'b000011111111;
20'b01011001110100011110: color_data = 12'b000011111111;
20'b01011001110100011111: color_data = 12'b000011111111;
20'b01011001110100100000: color_data = 12'b000011111111;
20'b01011010000011111010: color_data = 12'b000011111111;
20'b01011010000011111011: color_data = 12'b000011111111;
20'b01011010000011111100: color_data = 12'b000011111111;
20'b01011010000011111101: color_data = 12'b000011111111;
20'b01011010000011111110: color_data = 12'b000011111111;
20'b01011010000011111111: color_data = 12'b000011111111;
20'b01011010000100000000: color_data = 12'b000011111111;
20'b01011010000100000001: color_data = 12'b000011111111;
20'b01011010000100000010: color_data = 12'b000011111111;
20'b01011010000100000011: color_data = 12'b000011111111;
20'b01011010000100000100: color_data = 12'b000011111111;
20'b01011010000100000101: color_data = 12'b000011111111;
20'b01011010000100000110: color_data = 12'b000011111111;
20'b01011010000100000111: color_data = 12'b000011111111;
20'b01011010000100001000: color_data = 12'b000011111111;
20'b01011010000100001001: color_data = 12'b000011111111;
20'b01011010000100001010: color_data = 12'b000011111111;
20'b01011010000100001011: color_data = 12'b000011111111;
20'b01011010000100001111: color_data = 12'b000011111111;
20'b01011010000100010000: color_data = 12'b000011111111;
20'b01011010000100010001: color_data = 12'b000011111111;
20'b01011010000100010010: color_data = 12'b000011111111;
20'b01011010000100010011: color_data = 12'b000011111111;
20'b01011010000100010100: color_data = 12'b000011111111;
20'b01011010000100010101: color_data = 12'b000011111111;
20'b01011010000100010110: color_data = 12'b000011111111;
20'b01011010000100010111: color_data = 12'b000011111111;
20'b01011010000100011000: color_data = 12'b000011111111;
20'b01011010000100011001: color_data = 12'b000011111111;
20'b01011010000100011010: color_data = 12'b000011111111;
20'b01011010000100011011: color_data = 12'b000011111111;
20'b01011010000100011100: color_data = 12'b000011111111;
20'b01011010000100011101: color_data = 12'b000011111111;
20'b01011010000100011110: color_data = 12'b000011111111;
20'b01011010000100011111: color_data = 12'b000011111111;
20'b01011010000100100000: color_data = 12'b000011111111;
20'b01011010010011111010: color_data = 12'b000011111111;
20'b01011010010011111011: color_data = 12'b000011111111;
20'b01011010010011111100: color_data = 12'b000011111111;
20'b01011010010011111101: color_data = 12'b000011111111;
20'b01011010010011111110: color_data = 12'b000011111111;
20'b01011010010011111111: color_data = 12'b000011111111;
20'b01011010010100000000: color_data = 12'b000011111111;
20'b01011010010100000001: color_data = 12'b000011111111;
20'b01011010010100000010: color_data = 12'b000011111111;
20'b01011010010100000011: color_data = 12'b000011111111;
20'b01011010010100000100: color_data = 12'b000011111111;
20'b01011010010100000101: color_data = 12'b000011111111;
20'b01011010010100000110: color_data = 12'b000011111111;
20'b01011010010100000111: color_data = 12'b000011111111;
20'b01011010010100001000: color_data = 12'b000011111111;
20'b01011010010100001001: color_data = 12'b000011111111;
20'b01011010010100001010: color_data = 12'b000011111111;
20'b01011010010100001011: color_data = 12'b000011111111;
20'b01011010010100001111: color_data = 12'b000011111111;
20'b01011010010100010000: color_data = 12'b000011111111;
20'b01011010010100010001: color_data = 12'b000011111111;
20'b01011010010100010010: color_data = 12'b000011111111;
20'b01011010010100010011: color_data = 12'b000011111111;
20'b01011010010100010100: color_data = 12'b000011111111;
20'b01011010010100010101: color_data = 12'b000011111111;
20'b01011010010100010110: color_data = 12'b000011111111;
20'b01011010010100010111: color_data = 12'b000011111111;
20'b01011010010100011000: color_data = 12'b000011111111;
20'b01011010010100011001: color_data = 12'b000011111111;
20'b01011010010100011010: color_data = 12'b000011111111;
20'b01011010010100011011: color_data = 12'b000011111111;
20'b01011010010100011100: color_data = 12'b000011111111;
20'b01011010010100011101: color_data = 12'b000011111111;
20'b01011010010100011110: color_data = 12'b000011111111;
20'b01011010010100011111: color_data = 12'b000011111111;
20'b01011010010100100000: color_data = 12'b000011111111;
20'b01011010100011111010: color_data = 12'b000011111111;
20'b01011010100011111011: color_data = 12'b000011111111;
20'b01011010100011111100: color_data = 12'b000011111111;
20'b01011010100011111101: color_data = 12'b000011111111;
20'b01011010100011111110: color_data = 12'b000011111111;
20'b01011010100011111111: color_data = 12'b000011111111;
20'b01011010100100000000: color_data = 12'b000011111111;
20'b01011010100100000001: color_data = 12'b000011111111;
20'b01011010100100000010: color_data = 12'b000011111111;
20'b01011010100100000011: color_data = 12'b000011111111;
20'b01011010100100000100: color_data = 12'b000011111111;
20'b01011010100100000101: color_data = 12'b000011111111;
20'b01011010100100000110: color_data = 12'b000011111111;
20'b01011010100100000111: color_data = 12'b000011111111;
20'b01011010100100001000: color_data = 12'b000011111111;
20'b01011010100100001001: color_data = 12'b000011111111;
20'b01011010100100001010: color_data = 12'b000011111111;
20'b01011010100100001011: color_data = 12'b000011111111;
20'b01011010100100001111: color_data = 12'b000011111111;
20'b01011010100100010000: color_data = 12'b000011111111;
20'b01011010100100010001: color_data = 12'b000011111111;
20'b01011010100100010010: color_data = 12'b000011111111;
20'b01011010100100010011: color_data = 12'b000011111111;
20'b01011010100100010100: color_data = 12'b000011111111;
20'b01011010100100010101: color_data = 12'b000011111111;
20'b01011010100100010110: color_data = 12'b000011111111;
20'b01011010100100010111: color_data = 12'b000011111111;
20'b01011010100100011000: color_data = 12'b000011111111;
20'b01011010100100011001: color_data = 12'b000011111111;
20'b01011010100100011010: color_data = 12'b000011111111;
20'b01011010100100011011: color_data = 12'b000011111111;
20'b01011010100100011100: color_data = 12'b000011111111;
20'b01011010100100011101: color_data = 12'b000011111111;
20'b01011010100100011110: color_data = 12'b000011111111;
20'b01011010100100011111: color_data = 12'b000011111111;
20'b01011010100100100000: color_data = 12'b000011111111;
20'b01011010110011111010: color_data = 12'b000011111111;
20'b01011010110011111011: color_data = 12'b000011111111;
20'b01011010110011111100: color_data = 12'b000011111111;
20'b01011010110011111101: color_data = 12'b000011111111;
20'b01011010110011111110: color_data = 12'b000011111111;
20'b01011010110011111111: color_data = 12'b000011111111;
20'b01011010110100000000: color_data = 12'b000011111111;
20'b01011010110100000001: color_data = 12'b000011111111;
20'b01011010110100000010: color_data = 12'b000011111111;
20'b01011010110100000011: color_data = 12'b000011111111;
20'b01011010110100000100: color_data = 12'b000011111111;
20'b01011010110100000101: color_data = 12'b000011111111;
20'b01011010110100000110: color_data = 12'b000011111111;
20'b01011010110100000111: color_data = 12'b000011111111;
20'b01011010110100001000: color_data = 12'b000011111111;
20'b01011010110100001001: color_data = 12'b000011111111;
20'b01011010110100001010: color_data = 12'b000011111111;
20'b01011010110100001011: color_data = 12'b000011111111;
20'b01011010110100001111: color_data = 12'b000011111111;
20'b01011010110100010000: color_data = 12'b000011111111;
20'b01011010110100010001: color_data = 12'b000011111111;
20'b01011010110100010010: color_data = 12'b000011111111;
20'b01011010110100010011: color_data = 12'b000011111111;
20'b01011010110100010100: color_data = 12'b000011111111;
20'b01011010110100010101: color_data = 12'b000011111111;
20'b01011010110100010110: color_data = 12'b000011111111;
20'b01011010110100010111: color_data = 12'b000011111111;
20'b01011010110100011000: color_data = 12'b000011111111;
20'b01011010110100011001: color_data = 12'b000011111111;
20'b01011010110100011010: color_data = 12'b000011111111;
20'b01011010110100011011: color_data = 12'b000011111111;
20'b01011010110100011100: color_data = 12'b000011111111;
20'b01011010110100011101: color_data = 12'b000011111111;
20'b01011010110100011110: color_data = 12'b000011111111;
20'b01011010110100011111: color_data = 12'b000011111111;
20'b01011010110100100000: color_data = 12'b000011111111;
20'b01011011000011111010: color_data = 12'b000011111111;
20'b01011011000011111011: color_data = 12'b000011111111;
20'b01011011000011111100: color_data = 12'b000011111111;
20'b01011011000011111101: color_data = 12'b000011111111;
20'b01011011000011111110: color_data = 12'b000011111111;
20'b01011011000011111111: color_data = 12'b000011111111;
20'b01011011000100000000: color_data = 12'b000011111111;
20'b01011011000100000001: color_data = 12'b000011111111;
20'b01011011000100000010: color_data = 12'b000011111111;
20'b01011011000100000011: color_data = 12'b000011111111;
20'b01011011000100000100: color_data = 12'b000011111111;
20'b01011011000100000101: color_data = 12'b000011111111;
20'b01011011000100000110: color_data = 12'b000011111111;
20'b01011011000100000111: color_data = 12'b000011111111;
20'b01011011000100001000: color_data = 12'b000011111111;
20'b01011011000100001001: color_data = 12'b000011111111;
20'b01011011000100001010: color_data = 12'b000011111111;
20'b01011011000100001011: color_data = 12'b000011111111;
20'b01011011000100001111: color_data = 12'b000011111111;
20'b01011011000100010000: color_data = 12'b000011111111;
20'b01011011000100010001: color_data = 12'b000011111111;
20'b01011011000100010010: color_data = 12'b000011111111;
20'b01011011000100010011: color_data = 12'b000011111111;
20'b01011011000100010100: color_data = 12'b000011111111;
20'b01011011000100010101: color_data = 12'b000011111111;
20'b01011011000100010110: color_data = 12'b000011111111;
20'b01011011000100010111: color_data = 12'b000011111111;
20'b01011011000100011000: color_data = 12'b000011111111;
20'b01011011000100011001: color_data = 12'b000011111111;
20'b01011011000100011010: color_data = 12'b000011111111;
20'b01011011000100011011: color_data = 12'b000011111111;
20'b01011011000100011100: color_data = 12'b000011111111;
20'b01011011000100011101: color_data = 12'b000011111111;
20'b01011011000100011110: color_data = 12'b000011111111;
20'b01011011000100011111: color_data = 12'b000011111111;
20'b01011011000100100000: color_data = 12'b000011111111;
20'b01011011010011111010: color_data = 12'b000011111111;
20'b01011011010011111011: color_data = 12'b000011111111;
20'b01011011010011111100: color_data = 12'b000011111111;
20'b01011011010011111101: color_data = 12'b000011111111;
20'b01011011010011111110: color_data = 12'b000011111111;
20'b01011011010011111111: color_data = 12'b000011111111;
20'b01011011010100000000: color_data = 12'b000011111111;
20'b01011011010100000001: color_data = 12'b000011111111;
20'b01011011010100000010: color_data = 12'b000011111111;
20'b01011011010100000011: color_data = 12'b000011111111;
20'b01011011010100000100: color_data = 12'b000011111111;
20'b01011011010100000101: color_data = 12'b000011111111;
20'b01011011010100000110: color_data = 12'b000011111111;
20'b01011011010100000111: color_data = 12'b000011111111;
20'b01011011010100001000: color_data = 12'b000011111111;
20'b01011011010100001001: color_data = 12'b000011111111;
20'b01011011010100001010: color_data = 12'b000011111111;
20'b01011011010100001011: color_data = 12'b000011111111;
20'b01011011010100001111: color_data = 12'b000011111111;
20'b01011011010100010000: color_data = 12'b000011111111;
20'b01011011010100010001: color_data = 12'b000011111111;
20'b01011011010100010010: color_data = 12'b000011111111;
20'b01011011010100010011: color_data = 12'b000011111111;
20'b01011011010100010100: color_data = 12'b000011111111;
20'b01011011010100010101: color_data = 12'b000011111111;
20'b01011011010100010110: color_data = 12'b000011111111;
20'b01011011010100010111: color_data = 12'b000011111111;
20'b01011011010100011000: color_data = 12'b000011111111;
20'b01011011010100011001: color_data = 12'b000011111111;
20'b01011011010100011010: color_data = 12'b000011111111;
20'b01011011010100011011: color_data = 12'b000011111111;
20'b01011011010100011100: color_data = 12'b000011111111;
20'b01011011010100011101: color_data = 12'b000011111111;
20'b01011011010100011110: color_data = 12'b000011111111;
20'b01011011010100011111: color_data = 12'b000011111111;
20'b01011011010100100000: color_data = 12'b000011111111;
20'b01011011100011111010: color_data = 12'b000011111111;
20'b01011011100011111011: color_data = 12'b000011111111;
20'b01011011100011111100: color_data = 12'b000011111111;
20'b01011011100011111101: color_data = 12'b000011111111;
20'b01011011100011111110: color_data = 12'b000011111111;
20'b01011011100011111111: color_data = 12'b000011111111;
20'b01011011100100000000: color_data = 12'b000011111111;
20'b01011011100100000001: color_data = 12'b000011111111;
20'b01011011100100000010: color_data = 12'b000011111111;
20'b01011011100100000011: color_data = 12'b000011111111;
20'b01011011100100000100: color_data = 12'b000011111111;
20'b01011011100100000101: color_data = 12'b000011111111;
20'b01011011100100000110: color_data = 12'b000011111111;
20'b01011011100100000111: color_data = 12'b000011111111;
20'b01011011100100001000: color_data = 12'b000011111111;
20'b01011011100100001001: color_data = 12'b000011111111;
20'b01011011100100001010: color_data = 12'b000011111111;
20'b01011011100100001011: color_data = 12'b000011111111;
20'b01011011100100001111: color_data = 12'b000011111111;
20'b01011011100100010000: color_data = 12'b000011111111;
20'b01011011100100010001: color_data = 12'b000011111111;
20'b01011011100100010010: color_data = 12'b000011111111;
20'b01011011100100010011: color_data = 12'b000011111111;
20'b01011011100100010100: color_data = 12'b000011111111;
20'b01011011100100010101: color_data = 12'b000011111111;
20'b01011011100100010110: color_data = 12'b000011111111;
20'b01011011100100010111: color_data = 12'b000011111111;
20'b01011011100100011000: color_data = 12'b000011111111;
20'b01011011100100011001: color_data = 12'b000011111111;
20'b01011011100100011010: color_data = 12'b000011111111;
20'b01011011100100011011: color_data = 12'b000011111111;
20'b01011011100100011100: color_data = 12'b000011111111;
20'b01011011100100011101: color_data = 12'b000011111111;
20'b01011011100100011110: color_data = 12'b000011111111;
20'b01011011100100011111: color_data = 12'b000011111111;
20'b01011011100100100000: color_data = 12'b000011111111;
20'b01011011110011111010: color_data = 12'b000011111111;
20'b01011011110011111011: color_data = 12'b000011111111;
20'b01011011110011111100: color_data = 12'b000011111111;
20'b01011011110011111101: color_data = 12'b000011111111;
20'b01011011110011111110: color_data = 12'b000011111111;
20'b01011011110011111111: color_data = 12'b000011111111;
20'b01011011110100000000: color_data = 12'b000011111111;
20'b01011011110100000001: color_data = 12'b000011111111;
20'b01011011110100000010: color_data = 12'b000011111111;
20'b01011011110100000011: color_data = 12'b000011111111;
20'b01011011110100000100: color_data = 12'b000011111111;
20'b01011011110100000101: color_data = 12'b000011111111;
20'b01011011110100000110: color_data = 12'b000011111111;
20'b01011011110100000111: color_data = 12'b000011111111;
20'b01011011110100001000: color_data = 12'b000011111111;
20'b01011011110100001001: color_data = 12'b000011111111;
20'b01011011110100001010: color_data = 12'b000011111111;
20'b01011011110100001011: color_data = 12'b000011111111;
20'b01011011110100001111: color_data = 12'b000011111111;
20'b01011011110100010000: color_data = 12'b000011111111;
20'b01011011110100010001: color_data = 12'b000011111111;
20'b01011011110100010010: color_data = 12'b000011111111;
20'b01011011110100010011: color_data = 12'b000011111111;
20'b01011011110100010100: color_data = 12'b000011111111;
20'b01011011110100010101: color_data = 12'b000011111111;
20'b01011011110100010110: color_data = 12'b000011111111;
20'b01011011110100010111: color_data = 12'b000011111111;
20'b01011011110100011000: color_data = 12'b000011111111;
20'b01011011110100011001: color_data = 12'b000011111111;
20'b01011011110100011010: color_data = 12'b000011111111;
20'b01011011110100011011: color_data = 12'b000011111111;
20'b01011011110100011100: color_data = 12'b000011111111;
20'b01011011110100011101: color_data = 12'b000011111111;
20'b01011011110100011110: color_data = 12'b000011111111;
20'b01011011110100011111: color_data = 12'b000011111111;
20'b01011011110100100000: color_data = 12'b000011111111;
20'b01011100000011111010: color_data = 12'b000011111111;
20'b01011100000011111011: color_data = 12'b000011111111;
20'b01011100000011111100: color_data = 12'b000011111111;
20'b01011100000011111101: color_data = 12'b000011111111;
20'b01011100000011111110: color_data = 12'b000011111111;
20'b01011100000011111111: color_data = 12'b000011111111;
20'b01011100000100000000: color_data = 12'b000011111111;
20'b01011100000100000001: color_data = 12'b000011111111;
20'b01011100000100000010: color_data = 12'b000011111111;
20'b01011100000100000011: color_data = 12'b000011111111;
20'b01011100000100000100: color_data = 12'b000011111111;
20'b01011100000100000101: color_data = 12'b000011111111;
20'b01011100000100000110: color_data = 12'b000011111111;
20'b01011100000100000111: color_data = 12'b000011111111;
20'b01011100000100001000: color_data = 12'b000011111111;
20'b01011100000100001001: color_data = 12'b000011111111;
20'b01011100000100001010: color_data = 12'b000011111111;
20'b01011100000100001011: color_data = 12'b000011111111;
20'b01011100000100001111: color_data = 12'b000011111111;
20'b01011100000100010000: color_data = 12'b000011111111;
20'b01011100000100010001: color_data = 12'b000011111111;
20'b01011100000100010010: color_data = 12'b000011111111;
20'b01011100000100010011: color_data = 12'b000011111111;
20'b01011100000100010100: color_data = 12'b000011111111;
20'b01011100000100010101: color_data = 12'b000011111111;
20'b01011100000100010110: color_data = 12'b000011111111;
20'b01011100000100010111: color_data = 12'b000011111111;
20'b01011100000100011000: color_data = 12'b000011111111;
20'b01011100000100011001: color_data = 12'b000011111111;
20'b01011100000100011010: color_data = 12'b000011111111;
20'b01011100000100011011: color_data = 12'b000011111111;
20'b01011100000100011100: color_data = 12'b000011111111;
20'b01011100000100011101: color_data = 12'b000011111111;
20'b01011100000100011110: color_data = 12'b000011111111;
20'b01011100000100011111: color_data = 12'b000011111111;
20'b01011100000100100000: color_data = 12'b000011111111;
20'b01011100010011111010: color_data = 12'b000011111111;
20'b01011100010011111011: color_data = 12'b000011111111;
20'b01011100010011111100: color_data = 12'b000011111111;
20'b01011100010011111101: color_data = 12'b000011111111;
20'b01011100010011111110: color_data = 12'b000011111111;
20'b01011100010011111111: color_data = 12'b000011111111;
20'b01011100010100000000: color_data = 12'b000011111111;
20'b01011100010100000001: color_data = 12'b000011111111;
20'b01011100010100000010: color_data = 12'b000011111111;
20'b01011100010100000011: color_data = 12'b000011111111;
20'b01011100010100000100: color_data = 12'b000011111111;
20'b01011100010100000101: color_data = 12'b000011111111;
20'b01011100010100000110: color_data = 12'b000011111111;
20'b01011100010100000111: color_data = 12'b000011111111;
20'b01011100010100001000: color_data = 12'b000011111111;
20'b01011100010100001001: color_data = 12'b000011111111;
20'b01011100010100001010: color_data = 12'b000011111111;
20'b01011100010100001011: color_data = 12'b000011111111;
20'b01011100010100001111: color_data = 12'b000011111111;
20'b01011100010100010000: color_data = 12'b000011111111;
20'b01011100010100010001: color_data = 12'b000011111111;
20'b01011100010100010010: color_data = 12'b000011111111;
20'b01011100010100010011: color_data = 12'b000011111111;
20'b01011100010100010100: color_data = 12'b000011111111;
20'b01011100010100010101: color_data = 12'b000011111111;
20'b01011100010100010110: color_data = 12'b000011111111;
20'b01011100010100010111: color_data = 12'b000011111111;
20'b01011100010100011000: color_data = 12'b000011111111;
20'b01011100010100011001: color_data = 12'b000011111111;
20'b01011100010100011010: color_data = 12'b000011111111;
20'b01011100010100011011: color_data = 12'b000011111111;
20'b01011100010100011100: color_data = 12'b000011111111;
20'b01011100010100011101: color_data = 12'b000011111111;
20'b01011100010100011110: color_data = 12'b000011111111;
20'b01011100010100011111: color_data = 12'b000011111111;
20'b01011100010100100000: color_data = 12'b000011111111;
20'b01011100100011111010: color_data = 12'b000011111111;
20'b01011100100011111011: color_data = 12'b000011111111;
20'b01011100100011111100: color_data = 12'b000011111111;
20'b01011100100011111101: color_data = 12'b000011111111;
20'b01011100100011111110: color_data = 12'b000011111111;
20'b01011100100011111111: color_data = 12'b000011111111;
20'b01011100100100000000: color_data = 12'b000011111111;
20'b01011100100100000001: color_data = 12'b000011111111;
20'b01011100100100000010: color_data = 12'b000011111111;
20'b01011100100100000011: color_data = 12'b000011111111;
20'b01011100100100000100: color_data = 12'b000011111111;
20'b01011100100100000101: color_data = 12'b000011111111;
20'b01011100100100000110: color_data = 12'b000011111111;
20'b01011100100100000111: color_data = 12'b000011111111;
20'b01011100100100001000: color_data = 12'b000011111111;
20'b01011100100100001001: color_data = 12'b000011111111;
20'b01011100100100001010: color_data = 12'b000011111111;
20'b01011100100100001011: color_data = 12'b000011111111;
20'b01011100100100001111: color_data = 12'b000011111111;
20'b01011100100100010000: color_data = 12'b000011111111;
20'b01011100100100010001: color_data = 12'b000011111111;
20'b01011100100100010010: color_data = 12'b000011111111;
20'b01011100100100010011: color_data = 12'b000011111111;
20'b01011100100100010100: color_data = 12'b000011111111;
20'b01011100100100010101: color_data = 12'b000011111111;
20'b01011100100100010110: color_data = 12'b000011111111;
20'b01011100100100010111: color_data = 12'b000011111111;
20'b01011100100100011000: color_data = 12'b000011111111;
20'b01011100100100011001: color_data = 12'b000011111111;
20'b01011100100100011010: color_data = 12'b000011111111;
20'b01011100100100011011: color_data = 12'b000011111111;
20'b01011100100100011100: color_data = 12'b000011111111;
20'b01011100100100011101: color_data = 12'b000011111111;
20'b01011100100100011110: color_data = 12'b000011111111;
20'b01011100100100011111: color_data = 12'b000011111111;
20'b01011100100100100000: color_data = 12'b000011111111;
20'b01011100110011111010: color_data = 12'b000011111111;
20'b01011100110011111011: color_data = 12'b000011111111;
20'b01011100110011111100: color_data = 12'b000011111111;
20'b01011100110011111101: color_data = 12'b000011111111;
20'b01011100110011111110: color_data = 12'b000011111111;
20'b01011100110011111111: color_data = 12'b000011111111;
20'b01011100110100000000: color_data = 12'b000011111111;
20'b01011100110100000001: color_data = 12'b000011111111;
20'b01011100110100000010: color_data = 12'b000011111111;
20'b01011100110100000011: color_data = 12'b000011111111;
20'b01011100110100000100: color_data = 12'b000011111111;
20'b01011100110100000101: color_data = 12'b000011111111;
20'b01011100110100000110: color_data = 12'b000011111111;
20'b01011100110100000111: color_data = 12'b000011111111;
20'b01011100110100001000: color_data = 12'b000011111111;
20'b01011100110100001001: color_data = 12'b000011111111;
20'b01011100110100001010: color_data = 12'b000011111111;
20'b01011100110100001011: color_data = 12'b000011111111;
20'b01011100110100001111: color_data = 12'b000011111111;
20'b01011100110100010000: color_data = 12'b000011111111;
20'b01011100110100010001: color_data = 12'b000011111111;
20'b01011100110100010010: color_data = 12'b000011111111;
20'b01011100110100010011: color_data = 12'b000011111111;
20'b01011100110100010100: color_data = 12'b000011111111;
20'b01011100110100010101: color_data = 12'b000011111111;
20'b01011100110100010110: color_data = 12'b000011111111;
20'b01011100110100010111: color_data = 12'b000011111111;
20'b01011100110100011000: color_data = 12'b000011111111;
20'b01011100110100011001: color_data = 12'b000011111111;
20'b01011100110100011010: color_data = 12'b000011111111;
20'b01011100110100011011: color_data = 12'b000011111111;
20'b01011100110100011100: color_data = 12'b000011111111;
20'b01011100110100011101: color_data = 12'b000011111111;
20'b01011100110100011110: color_data = 12'b000011111111;
20'b01011100110100011111: color_data = 12'b000011111111;
20'b01011100110100100000: color_data = 12'b000011111111;
20'b01011101000011111010: color_data = 12'b000011111111;
20'b01011101000011111011: color_data = 12'b000011111111;
20'b01011101000011111100: color_data = 12'b000011111111;
20'b01011101000011111101: color_data = 12'b000011111111;
20'b01011101000011111110: color_data = 12'b000011111111;
20'b01011101000011111111: color_data = 12'b000011111111;
20'b01011101000100000000: color_data = 12'b000011111111;
20'b01011101000100000001: color_data = 12'b000011111111;
20'b01011101000100000010: color_data = 12'b000011111111;
20'b01011101000100000011: color_data = 12'b000011111111;
20'b01011101000100000100: color_data = 12'b000011111111;
20'b01011101000100000101: color_data = 12'b000011111111;
20'b01011101000100000110: color_data = 12'b000011111111;
20'b01011101000100000111: color_data = 12'b000011111111;
20'b01011101000100001000: color_data = 12'b000011111111;
20'b01011101000100001001: color_data = 12'b000011111111;
20'b01011101000100001010: color_data = 12'b000011111111;
20'b01011101000100001011: color_data = 12'b000011111111;
20'b01011101000100001111: color_data = 12'b000011111111;
20'b01011101000100010000: color_data = 12'b000011111111;
20'b01011101000100010001: color_data = 12'b000011111111;
20'b01011101000100010010: color_data = 12'b000011111111;
20'b01011101000100010011: color_data = 12'b000011111111;
20'b01011101000100010100: color_data = 12'b000011111111;
20'b01011101000100010101: color_data = 12'b000011111111;
20'b01011101000100010110: color_data = 12'b000011111111;
20'b01011101000100010111: color_data = 12'b000011111111;
20'b01011101000100011000: color_data = 12'b000011111111;
20'b01011101000100011001: color_data = 12'b000011111111;
20'b01011101000100011010: color_data = 12'b000011111111;
20'b01011101000100011011: color_data = 12'b000011111111;
20'b01011101000100011100: color_data = 12'b000011111111;
20'b01011101000100011101: color_data = 12'b000011111111;
20'b01011101000100011110: color_data = 12'b000011111111;
20'b01011101000100011111: color_data = 12'b000011111111;
20'b01011101000100100000: color_data = 12'b000011111111;
20'b01011101010011111010: color_data = 12'b000011111111;
20'b01011101010011111011: color_data = 12'b000011111111;
20'b01011101010011111100: color_data = 12'b000011111111;
20'b01011101010011111101: color_data = 12'b000011111111;
20'b01011101010011111110: color_data = 12'b000011111111;
20'b01011101010011111111: color_data = 12'b000011111111;
20'b01011101010100000000: color_data = 12'b000011111111;
20'b01011101010100000001: color_data = 12'b000011111111;
20'b01011101010100000010: color_data = 12'b000011111111;
20'b01011101010100000011: color_data = 12'b000011111111;
20'b01011101010100000100: color_data = 12'b000011111111;
20'b01011101010100000101: color_data = 12'b000011111111;
20'b01011101010100000110: color_data = 12'b000011111111;
20'b01011101010100000111: color_data = 12'b000011111111;
20'b01011101010100001000: color_data = 12'b000011111111;
20'b01011101010100001001: color_data = 12'b000011111111;
20'b01011101010100001010: color_data = 12'b000011111111;
20'b01011101010100001011: color_data = 12'b000011111111;
20'b01011101010100001111: color_data = 12'b000011111111;
20'b01011101010100010000: color_data = 12'b000011111111;
20'b01011101010100010001: color_data = 12'b000011111111;
20'b01011101010100010010: color_data = 12'b000011111111;
20'b01011101010100010011: color_data = 12'b000011111111;
20'b01011101010100010100: color_data = 12'b000011111111;
20'b01011101010100010101: color_data = 12'b000011111111;
20'b01011101010100010110: color_data = 12'b000011111111;
20'b01011101010100010111: color_data = 12'b000011111111;
20'b01011101010100011000: color_data = 12'b000011111111;
20'b01011101010100011001: color_data = 12'b000011111111;
20'b01011101010100011010: color_data = 12'b000011111111;
20'b01011101010100011011: color_data = 12'b000011111111;
20'b01011101010100011100: color_data = 12'b000011111111;
20'b01011101010100011101: color_data = 12'b000011111111;
20'b01011101010100011110: color_data = 12'b000011111111;
20'b01011101010100011111: color_data = 12'b000011111111;
20'b01011101010100100000: color_data = 12'b000011111111;
20'b01011101100011111010: color_data = 12'b000011111111;
20'b01011101100011111011: color_data = 12'b000011111111;
20'b01011101100011111100: color_data = 12'b000011111111;
20'b01011101100011111101: color_data = 12'b000011111111;
20'b01011101100011111110: color_data = 12'b000011111111;
20'b01011101100011111111: color_data = 12'b000011111111;
20'b01011101100100000000: color_data = 12'b000011111111;
20'b01011101100100000001: color_data = 12'b000011111111;
20'b01011101100100000010: color_data = 12'b000011111111;
20'b01011101100100000011: color_data = 12'b000011111111;
20'b01011101100100000100: color_data = 12'b000011111111;
20'b01011101100100000101: color_data = 12'b000011111111;
20'b01011101100100000110: color_data = 12'b000011111111;
20'b01011101100100000111: color_data = 12'b000011111111;
20'b01011101100100001000: color_data = 12'b000011111111;
20'b01011101100100001001: color_data = 12'b000011111111;
20'b01011101100100001010: color_data = 12'b000011111111;
20'b01011101100100001011: color_data = 12'b000011111111;
20'b01011101100100001111: color_data = 12'b000011111111;
20'b01011101100100010000: color_data = 12'b000011111111;
20'b01011101100100010001: color_data = 12'b000011111111;
20'b01011101100100010010: color_data = 12'b000011111111;
20'b01011101100100010011: color_data = 12'b000011111111;
20'b01011101100100010100: color_data = 12'b000011111111;
20'b01011101100100010101: color_data = 12'b000011111111;
20'b01011101100100010110: color_data = 12'b000011111111;
20'b01011101100100010111: color_data = 12'b000011111111;
20'b01011101100100011000: color_data = 12'b000011111111;
20'b01011101100100011001: color_data = 12'b000011111111;
20'b01011101100100011010: color_data = 12'b000011111111;
20'b01011101100100011011: color_data = 12'b000011111111;
20'b01011101100100011100: color_data = 12'b000011111111;
20'b01011101100100011101: color_data = 12'b000011111111;
20'b01011101100100011110: color_data = 12'b000011111111;
20'b01011101100100011111: color_data = 12'b000011111111;
20'b01011101100100100000: color_data = 12'b000011111111;
20'b01011101110011111010: color_data = 12'b000011111111;
20'b01011101110011111011: color_data = 12'b000011111111;
20'b01011101110011111100: color_data = 12'b000011111111;
20'b01011101110011111101: color_data = 12'b000011111111;
20'b01011101110011111110: color_data = 12'b000011111111;
20'b01011101110011111111: color_data = 12'b000011111111;
20'b01011101110100000000: color_data = 12'b000011111111;
20'b01011101110100000001: color_data = 12'b000011111111;
20'b01011101110100000010: color_data = 12'b000011111111;
20'b01011101110100000011: color_data = 12'b000011111111;
20'b01011101110100000100: color_data = 12'b000011111111;
20'b01011101110100000101: color_data = 12'b000011111111;
20'b01011101110100000110: color_data = 12'b000011111111;
20'b01011101110100000111: color_data = 12'b000011111111;
20'b01011101110100001000: color_data = 12'b000011111111;
20'b01011101110100001001: color_data = 12'b000011111111;
20'b01011101110100001010: color_data = 12'b000011111111;
20'b01011101110100001011: color_data = 12'b000011111111;
20'b01011101110100001111: color_data = 12'b000011111111;
20'b01011101110100010000: color_data = 12'b000011111111;
20'b01011101110100010001: color_data = 12'b000011111111;
20'b01011101110100010010: color_data = 12'b000011111111;
20'b01011101110100010011: color_data = 12'b000011111111;
20'b01011101110100010100: color_data = 12'b000011111111;
20'b01011101110100010101: color_data = 12'b000011111111;
20'b01011101110100010110: color_data = 12'b000011111111;
20'b01011101110100010111: color_data = 12'b000011111111;
20'b01011101110100011000: color_data = 12'b000011111111;
20'b01011101110100011001: color_data = 12'b000011111111;
20'b01011101110100011010: color_data = 12'b000011111111;
20'b01011101110100011011: color_data = 12'b000011111111;
20'b01011101110100011100: color_data = 12'b000011111111;
20'b01011101110100011101: color_data = 12'b000011111111;
20'b01011101110100011110: color_data = 12'b000011111111;
20'b01011101110100011111: color_data = 12'b000011111111;
20'b01011101110100100000: color_data = 12'b000011111111;
20'b01011110110011111010: color_data = 12'b000011111111;
20'b01011110110011111011: color_data = 12'b000011111111;
20'b01011110110011111100: color_data = 12'b000011111111;
20'b01011110110011111101: color_data = 12'b000011111111;
20'b01011110110011111110: color_data = 12'b000011111111;
20'b01011110110011111111: color_data = 12'b000011111111;
20'b01011110110100000000: color_data = 12'b000011111111;
20'b01011110110100000001: color_data = 12'b000011111111;
20'b01011110110100000010: color_data = 12'b000011111111;
20'b01011110110100000011: color_data = 12'b000011111111;
20'b01011110110100000100: color_data = 12'b000011111111;
20'b01011110110100000101: color_data = 12'b000011111111;
20'b01011110110100000110: color_data = 12'b000011111111;
20'b01011110110100000111: color_data = 12'b000011111111;
20'b01011110110100001000: color_data = 12'b000011111111;
20'b01011110110100001001: color_data = 12'b000011111111;
20'b01011110110100001010: color_data = 12'b000011111111;
20'b01011110110100001011: color_data = 12'b000011111111;
20'b01011110110100001111: color_data = 12'b000011111111;
20'b01011110110100010000: color_data = 12'b000011111111;
20'b01011110110100010001: color_data = 12'b000011111111;
20'b01011110110100010010: color_data = 12'b000011111111;
20'b01011110110100010011: color_data = 12'b000011111111;
20'b01011110110100010100: color_data = 12'b000011111111;
20'b01011110110100010101: color_data = 12'b000011111111;
20'b01011110110100010110: color_data = 12'b000011111111;
20'b01011110110100010111: color_data = 12'b000011111111;
20'b01011110110100011000: color_data = 12'b000011111111;
20'b01011110110100011001: color_data = 12'b000011111111;
20'b01011110110100011010: color_data = 12'b000011111111;
20'b01011110110100011011: color_data = 12'b000011111111;
20'b01011110110100011100: color_data = 12'b000011111111;
20'b01011110110100011101: color_data = 12'b000011111111;
20'b01011110110100011110: color_data = 12'b000011111111;
20'b01011110110100011111: color_data = 12'b000011111111;
20'b01011110110100100000: color_data = 12'b000011111111;
20'b01011110110100100100: color_data = 12'b000001101111;
20'b01011110110100100101: color_data = 12'b000001101111;
20'b01011110110100100110: color_data = 12'b000001101111;
20'b01011110110100100111: color_data = 12'b000001101111;
20'b01011110110100101000: color_data = 12'b000001101111;
20'b01011110110100101001: color_data = 12'b000001101111;
20'b01011110110100101010: color_data = 12'b000001101111;
20'b01011110110100101011: color_data = 12'b000001101111;
20'b01011110110100101100: color_data = 12'b000001101111;
20'b01011110110100101101: color_data = 12'b000001101111;
20'b01011110110100101110: color_data = 12'b000001101111;
20'b01011110110100101111: color_data = 12'b000001101111;
20'b01011110110100110000: color_data = 12'b000001101111;
20'b01011110110100110001: color_data = 12'b000001101111;
20'b01011110110100110010: color_data = 12'b000001101111;
20'b01011110110100110011: color_data = 12'b000001101111;
20'b01011110110100110100: color_data = 12'b000001101111;
20'b01011110110100110101: color_data = 12'b000001101111;
20'b01011110110100111001: color_data = 12'b000011110000;
20'b01011110110100111010: color_data = 12'b000011110000;
20'b01011110110100111011: color_data = 12'b000011110000;
20'b01011110110100111100: color_data = 12'b000011110000;
20'b01011110110100111101: color_data = 12'b000011110000;
20'b01011110110100111110: color_data = 12'b000011110000;
20'b01011110110100111111: color_data = 12'b000011110000;
20'b01011110110101000000: color_data = 12'b000011110000;
20'b01011110110101000001: color_data = 12'b000011110000;
20'b01011110110101000010: color_data = 12'b000011110000;
20'b01011110110101000011: color_data = 12'b000011110000;
20'b01011110110101000100: color_data = 12'b000011110000;
20'b01011110110101000101: color_data = 12'b000011110000;
20'b01011110110101000110: color_data = 12'b000011110000;
20'b01011110110101000111: color_data = 12'b000011110000;
20'b01011110110101001000: color_data = 12'b000011110000;
20'b01011110110101001001: color_data = 12'b000011110000;
20'b01011110110101001010: color_data = 12'b000011110000;
20'b01011110110101100011: color_data = 12'b111100001111;
20'b01011110110101100100: color_data = 12'b111100001111;
20'b01011110110101100101: color_data = 12'b111100001111;
20'b01011110110101100110: color_data = 12'b111100001111;
20'b01011110110101100111: color_data = 12'b111100001111;
20'b01011110110101101000: color_data = 12'b111100001111;
20'b01011110110101101001: color_data = 12'b111100001111;
20'b01011110110101101010: color_data = 12'b111100001111;
20'b01011110110101101011: color_data = 12'b111100001111;
20'b01011110110101101100: color_data = 12'b111100001111;
20'b01011110110101101101: color_data = 12'b111100001111;
20'b01011110110101101110: color_data = 12'b111100001111;
20'b01011110110101101111: color_data = 12'b111100001111;
20'b01011110110101110000: color_data = 12'b111100001111;
20'b01011110110101110001: color_data = 12'b111100001111;
20'b01011110110101110010: color_data = 12'b111100001111;
20'b01011110110101110011: color_data = 12'b111100001111;
20'b01011110110101110100: color_data = 12'b111100001111;
20'b01011110110110001101: color_data = 12'b111100000000;
20'b01011110110110001110: color_data = 12'b111100000000;
20'b01011110110110001111: color_data = 12'b111100000000;
20'b01011110110110010000: color_data = 12'b111100000000;
20'b01011110110110010001: color_data = 12'b111100000000;
20'b01011110110110010010: color_data = 12'b111100000000;
20'b01011110110110010011: color_data = 12'b111100000000;
20'b01011110110110010100: color_data = 12'b111100000000;
20'b01011110110110010101: color_data = 12'b111100000000;
20'b01011110110110010110: color_data = 12'b111100000000;
20'b01011110110110010111: color_data = 12'b111100000000;
20'b01011110110110011000: color_data = 12'b111100000000;
20'b01011110110110011001: color_data = 12'b111100000000;
20'b01011110110110011010: color_data = 12'b111100000000;
20'b01011110110110011011: color_data = 12'b111100000000;
20'b01011110110110011100: color_data = 12'b111100000000;
20'b01011110110110011101: color_data = 12'b111100000000;
20'b01011110110110011110: color_data = 12'b111100000000;
20'b01011111000011111010: color_data = 12'b000011111111;
20'b01011111000011111011: color_data = 12'b000011111111;
20'b01011111000011111100: color_data = 12'b000011111111;
20'b01011111000011111101: color_data = 12'b000011111111;
20'b01011111000011111110: color_data = 12'b000011111111;
20'b01011111000011111111: color_data = 12'b000011111111;
20'b01011111000100000000: color_data = 12'b000011111111;
20'b01011111000100000001: color_data = 12'b000011111111;
20'b01011111000100000010: color_data = 12'b000011111111;
20'b01011111000100000011: color_data = 12'b000011111111;
20'b01011111000100000100: color_data = 12'b000011111111;
20'b01011111000100000101: color_data = 12'b000011111111;
20'b01011111000100000110: color_data = 12'b000011111111;
20'b01011111000100000111: color_data = 12'b000011111111;
20'b01011111000100001000: color_data = 12'b000011111111;
20'b01011111000100001001: color_data = 12'b000011111111;
20'b01011111000100001010: color_data = 12'b000011111111;
20'b01011111000100001011: color_data = 12'b000011111111;
20'b01011111000100001111: color_data = 12'b000011111111;
20'b01011111000100010000: color_data = 12'b000011111111;
20'b01011111000100010001: color_data = 12'b000011111111;
20'b01011111000100010010: color_data = 12'b000011111111;
20'b01011111000100010011: color_data = 12'b000011111111;
20'b01011111000100010100: color_data = 12'b000011111111;
20'b01011111000100010101: color_data = 12'b000011111111;
20'b01011111000100010110: color_data = 12'b000011111111;
20'b01011111000100010111: color_data = 12'b000011111111;
20'b01011111000100011000: color_data = 12'b000011111111;
20'b01011111000100011001: color_data = 12'b000011111111;
20'b01011111000100011010: color_data = 12'b000011111111;
20'b01011111000100011011: color_data = 12'b000011111111;
20'b01011111000100011100: color_data = 12'b000011111111;
20'b01011111000100011101: color_data = 12'b000011111111;
20'b01011111000100011110: color_data = 12'b000011111111;
20'b01011111000100011111: color_data = 12'b000011111111;
20'b01011111000100100000: color_data = 12'b000011111111;
20'b01011111000100100100: color_data = 12'b000001101111;
20'b01011111000100100101: color_data = 12'b000001101111;
20'b01011111000100100110: color_data = 12'b000001101111;
20'b01011111000100100111: color_data = 12'b000001101111;
20'b01011111000100101000: color_data = 12'b000001101111;
20'b01011111000100101001: color_data = 12'b000001101111;
20'b01011111000100101010: color_data = 12'b000001101111;
20'b01011111000100101011: color_data = 12'b000001101111;
20'b01011111000100101100: color_data = 12'b000001101111;
20'b01011111000100101101: color_data = 12'b000001101111;
20'b01011111000100101110: color_data = 12'b000001101111;
20'b01011111000100101111: color_data = 12'b000001101111;
20'b01011111000100110000: color_data = 12'b000001101111;
20'b01011111000100110001: color_data = 12'b000001101111;
20'b01011111000100110010: color_data = 12'b000001101111;
20'b01011111000100110011: color_data = 12'b000001101111;
20'b01011111000100110100: color_data = 12'b000001101111;
20'b01011111000100110101: color_data = 12'b000001101111;
20'b01011111000100111001: color_data = 12'b000011110000;
20'b01011111000100111010: color_data = 12'b000011110000;
20'b01011111000100111011: color_data = 12'b000011110000;
20'b01011111000100111100: color_data = 12'b000011110000;
20'b01011111000100111101: color_data = 12'b000011110000;
20'b01011111000100111110: color_data = 12'b000011110000;
20'b01011111000100111111: color_data = 12'b000011110000;
20'b01011111000101000000: color_data = 12'b000011110000;
20'b01011111000101000001: color_data = 12'b000011110000;
20'b01011111000101000010: color_data = 12'b000011110000;
20'b01011111000101000011: color_data = 12'b000011110000;
20'b01011111000101000100: color_data = 12'b000011110000;
20'b01011111000101000101: color_data = 12'b000011110000;
20'b01011111000101000110: color_data = 12'b000011110000;
20'b01011111000101000111: color_data = 12'b000011110000;
20'b01011111000101001000: color_data = 12'b000011110000;
20'b01011111000101001001: color_data = 12'b000011110000;
20'b01011111000101001010: color_data = 12'b000011110000;
20'b01011111000101100011: color_data = 12'b111100001111;
20'b01011111000101100100: color_data = 12'b111100001111;
20'b01011111000101100101: color_data = 12'b111100001111;
20'b01011111000101100110: color_data = 12'b111100001111;
20'b01011111000101100111: color_data = 12'b111100001111;
20'b01011111000101101000: color_data = 12'b111100001111;
20'b01011111000101101001: color_data = 12'b111100001111;
20'b01011111000101101010: color_data = 12'b111100001111;
20'b01011111000101101011: color_data = 12'b111100001111;
20'b01011111000101101100: color_data = 12'b111100001111;
20'b01011111000101101101: color_data = 12'b111100001111;
20'b01011111000101101110: color_data = 12'b111100001111;
20'b01011111000101101111: color_data = 12'b111100001111;
20'b01011111000101110000: color_data = 12'b111100001111;
20'b01011111000101110001: color_data = 12'b111100001111;
20'b01011111000101110010: color_data = 12'b111100001111;
20'b01011111000101110011: color_data = 12'b111100001111;
20'b01011111000101110100: color_data = 12'b111100001111;
20'b01011111000110001101: color_data = 12'b111100000000;
20'b01011111000110001110: color_data = 12'b111100000000;
20'b01011111000110001111: color_data = 12'b111100000000;
20'b01011111000110010000: color_data = 12'b111100000000;
20'b01011111000110010001: color_data = 12'b111100000000;
20'b01011111000110010010: color_data = 12'b111100000000;
20'b01011111000110010011: color_data = 12'b111100000000;
20'b01011111000110010100: color_data = 12'b111100000000;
20'b01011111000110010101: color_data = 12'b111100000000;
20'b01011111000110010110: color_data = 12'b111100000000;
20'b01011111000110010111: color_data = 12'b111100000000;
20'b01011111000110011000: color_data = 12'b111100000000;
20'b01011111000110011001: color_data = 12'b111100000000;
20'b01011111000110011010: color_data = 12'b111100000000;
20'b01011111000110011011: color_data = 12'b111100000000;
20'b01011111000110011100: color_data = 12'b111100000000;
20'b01011111000110011101: color_data = 12'b111100000000;
20'b01011111000110011110: color_data = 12'b111100000000;
20'b01011111010011111010: color_data = 12'b000011111111;
20'b01011111010011111011: color_data = 12'b000011111111;
20'b01011111010011111100: color_data = 12'b000011111111;
20'b01011111010011111101: color_data = 12'b000011111111;
20'b01011111010011111110: color_data = 12'b000011111111;
20'b01011111010011111111: color_data = 12'b000011111111;
20'b01011111010100000000: color_data = 12'b000011111111;
20'b01011111010100000001: color_data = 12'b000011111111;
20'b01011111010100000010: color_data = 12'b000011111111;
20'b01011111010100000011: color_data = 12'b000011111111;
20'b01011111010100000100: color_data = 12'b000011111111;
20'b01011111010100000101: color_data = 12'b000011111111;
20'b01011111010100000110: color_data = 12'b000011111111;
20'b01011111010100000111: color_data = 12'b000011111111;
20'b01011111010100001000: color_data = 12'b000011111111;
20'b01011111010100001001: color_data = 12'b000011111111;
20'b01011111010100001010: color_data = 12'b000011111111;
20'b01011111010100001011: color_data = 12'b000011111111;
20'b01011111010100001111: color_data = 12'b000011111111;
20'b01011111010100010000: color_data = 12'b000011111111;
20'b01011111010100010001: color_data = 12'b000011111111;
20'b01011111010100010010: color_data = 12'b000011111111;
20'b01011111010100010011: color_data = 12'b000011111111;
20'b01011111010100010100: color_data = 12'b000011111111;
20'b01011111010100010101: color_data = 12'b000011111111;
20'b01011111010100010110: color_data = 12'b000011111111;
20'b01011111010100010111: color_data = 12'b000011111111;
20'b01011111010100011000: color_data = 12'b000011111111;
20'b01011111010100011001: color_data = 12'b000011111111;
20'b01011111010100011010: color_data = 12'b000011111111;
20'b01011111010100011011: color_data = 12'b000011111111;
20'b01011111010100011100: color_data = 12'b000011111111;
20'b01011111010100011101: color_data = 12'b000011111111;
20'b01011111010100011110: color_data = 12'b000011111111;
20'b01011111010100011111: color_data = 12'b000011111111;
20'b01011111010100100000: color_data = 12'b000011111111;
20'b01011111010100100100: color_data = 12'b000001101111;
20'b01011111010100100101: color_data = 12'b000001101111;
20'b01011111010100100110: color_data = 12'b000001101111;
20'b01011111010100100111: color_data = 12'b000001101111;
20'b01011111010100101000: color_data = 12'b000001101111;
20'b01011111010100101001: color_data = 12'b000001101111;
20'b01011111010100101010: color_data = 12'b000001101111;
20'b01011111010100101011: color_data = 12'b000001101111;
20'b01011111010100101100: color_data = 12'b000001101111;
20'b01011111010100101101: color_data = 12'b000001101111;
20'b01011111010100101110: color_data = 12'b000001101111;
20'b01011111010100101111: color_data = 12'b000001101111;
20'b01011111010100110000: color_data = 12'b000001101111;
20'b01011111010100110001: color_data = 12'b000001101111;
20'b01011111010100110010: color_data = 12'b000001101111;
20'b01011111010100110011: color_data = 12'b000001101111;
20'b01011111010100110100: color_data = 12'b000001101111;
20'b01011111010100110101: color_data = 12'b000001101111;
20'b01011111010100111001: color_data = 12'b000011110000;
20'b01011111010100111010: color_data = 12'b000011110000;
20'b01011111010100111011: color_data = 12'b000011110000;
20'b01011111010100111100: color_data = 12'b000011110000;
20'b01011111010100111101: color_data = 12'b000011110000;
20'b01011111010100111110: color_data = 12'b000011110000;
20'b01011111010100111111: color_data = 12'b000011110000;
20'b01011111010101000000: color_data = 12'b000011110000;
20'b01011111010101000001: color_data = 12'b000011110000;
20'b01011111010101000010: color_data = 12'b000011110000;
20'b01011111010101000011: color_data = 12'b000011110000;
20'b01011111010101000100: color_data = 12'b000011110000;
20'b01011111010101000101: color_data = 12'b000011110000;
20'b01011111010101000110: color_data = 12'b000011110000;
20'b01011111010101000111: color_data = 12'b000011110000;
20'b01011111010101001000: color_data = 12'b000011110000;
20'b01011111010101001001: color_data = 12'b000011110000;
20'b01011111010101001010: color_data = 12'b000011110000;
20'b01011111010101100011: color_data = 12'b111100001111;
20'b01011111010101100100: color_data = 12'b111100001111;
20'b01011111010101100101: color_data = 12'b111100001111;
20'b01011111010101100110: color_data = 12'b111100001111;
20'b01011111010101100111: color_data = 12'b111100001111;
20'b01011111010101101000: color_data = 12'b111100001111;
20'b01011111010101101001: color_data = 12'b111100001111;
20'b01011111010101101010: color_data = 12'b111100001111;
20'b01011111010101101011: color_data = 12'b111100001111;
20'b01011111010101101100: color_data = 12'b111100001111;
20'b01011111010101101101: color_data = 12'b111100001111;
20'b01011111010101101110: color_data = 12'b111100001111;
20'b01011111010101101111: color_data = 12'b111100001111;
20'b01011111010101110000: color_data = 12'b111100001111;
20'b01011111010101110001: color_data = 12'b111100001111;
20'b01011111010101110010: color_data = 12'b111100001111;
20'b01011111010101110011: color_data = 12'b111100001111;
20'b01011111010101110100: color_data = 12'b111100001111;
20'b01011111010110001101: color_data = 12'b111100000000;
20'b01011111010110001110: color_data = 12'b111100000000;
20'b01011111010110001111: color_data = 12'b111100000000;
20'b01011111010110010000: color_data = 12'b111100000000;
20'b01011111010110010001: color_data = 12'b111100000000;
20'b01011111010110010010: color_data = 12'b111100000000;
20'b01011111010110010011: color_data = 12'b111100000000;
20'b01011111010110010100: color_data = 12'b111100000000;
20'b01011111010110010101: color_data = 12'b111100000000;
20'b01011111010110010110: color_data = 12'b111100000000;
20'b01011111010110010111: color_data = 12'b111100000000;
20'b01011111010110011000: color_data = 12'b111100000000;
20'b01011111010110011001: color_data = 12'b111100000000;
20'b01011111010110011010: color_data = 12'b111100000000;
20'b01011111010110011011: color_data = 12'b111100000000;
20'b01011111010110011100: color_data = 12'b111100000000;
20'b01011111010110011101: color_data = 12'b111100000000;
20'b01011111010110011110: color_data = 12'b111100000000;
20'b01011111100011111010: color_data = 12'b000011111111;
20'b01011111100011111011: color_data = 12'b000011111111;
20'b01011111100011111100: color_data = 12'b000011111111;
20'b01011111100011111101: color_data = 12'b000011111111;
20'b01011111100011111110: color_data = 12'b000011111111;
20'b01011111100011111111: color_data = 12'b000011111111;
20'b01011111100100000000: color_data = 12'b000011111111;
20'b01011111100100000001: color_data = 12'b000011111111;
20'b01011111100100000010: color_data = 12'b000011111111;
20'b01011111100100000011: color_data = 12'b000011111111;
20'b01011111100100000100: color_data = 12'b000011111111;
20'b01011111100100000101: color_data = 12'b000011111111;
20'b01011111100100000110: color_data = 12'b000011111111;
20'b01011111100100000111: color_data = 12'b000011111111;
20'b01011111100100001000: color_data = 12'b000011111111;
20'b01011111100100001001: color_data = 12'b000011111111;
20'b01011111100100001010: color_data = 12'b000011111111;
20'b01011111100100001011: color_data = 12'b000011111111;
20'b01011111100100001111: color_data = 12'b000011111111;
20'b01011111100100010000: color_data = 12'b000011111111;
20'b01011111100100010001: color_data = 12'b000011111111;
20'b01011111100100010010: color_data = 12'b000011111111;
20'b01011111100100010011: color_data = 12'b000011111111;
20'b01011111100100010100: color_data = 12'b000011111111;
20'b01011111100100010101: color_data = 12'b000011111111;
20'b01011111100100010110: color_data = 12'b000011111111;
20'b01011111100100010111: color_data = 12'b000011111111;
20'b01011111100100011000: color_data = 12'b000011111111;
20'b01011111100100011001: color_data = 12'b000011111111;
20'b01011111100100011010: color_data = 12'b000011111111;
20'b01011111100100011011: color_data = 12'b000011111111;
20'b01011111100100011100: color_data = 12'b000011111111;
20'b01011111100100011101: color_data = 12'b000011111111;
20'b01011111100100011110: color_data = 12'b000011111111;
20'b01011111100100011111: color_data = 12'b000011111111;
20'b01011111100100100000: color_data = 12'b000011111111;
20'b01011111100100100100: color_data = 12'b000001101111;
20'b01011111100100100101: color_data = 12'b000001101111;
20'b01011111100100100110: color_data = 12'b000001101111;
20'b01011111100100100111: color_data = 12'b000001101111;
20'b01011111100100101000: color_data = 12'b000001101111;
20'b01011111100100101001: color_data = 12'b000001101111;
20'b01011111100100101010: color_data = 12'b000001101111;
20'b01011111100100101011: color_data = 12'b000001101111;
20'b01011111100100101100: color_data = 12'b000001101111;
20'b01011111100100101101: color_data = 12'b000001101111;
20'b01011111100100101110: color_data = 12'b000001101111;
20'b01011111100100101111: color_data = 12'b000001101111;
20'b01011111100100110000: color_data = 12'b000001101111;
20'b01011111100100110001: color_data = 12'b000001101111;
20'b01011111100100110010: color_data = 12'b000001101111;
20'b01011111100100110011: color_data = 12'b000001101111;
20'b01011111100100110100: color_data = 12'b000001101111;
20'b01011111100100110101: color_data = 12'b000001101111;
20'b01011111100100111001: color_data = 12'b000011110000;
20'b01011111100100111010: color_data = 12'b000011110000;
20'b01011111100100111011: color_data = 12'b000011110000;
20'b01011111100100111100: color_data = 12'b000011110000;
20'b01011111100100111101: color_data = 12'b000011110000;
20'b01011111100100111110: color_data = 12'b000011110000;
20'b01011111100100111111: color_data = 12'b000011110000;
20'b01011111100101000000: color_data = 12'b000011110000;
20'b01011111100101000001: color_data = 12'b000011110000;
20'b01011111100101000010: color_data = 12'b000011110000;
20'b01011111100101000011: color_data = 12'b000011110000;
20'b01011111100101000100: color_data = 12'b000011110000;
20'b01011111100101000101: color_data = 12'b000011110000;
20'b01011111100101000110: color_data = 12'b000011110000;
20'b01011111100101000111: color_data = 12'b000011110000;
20'b01011111100101001000: color_data = 12'b000011110000;
20'b01011111100101001001: color_data = 12'b000011110000;
20'b01011111100101001010: color_data = 12'b000011110000;
20'b01011111100101100011: color_data = 12'b111100001111;
20'b01011111100101100100: color_data = 12'b111100001111;
20'b01011111100101100101: color_data = 12'b111100001111;
20'b01011111100101100110: color_data = 12'b111100001111;
20'b01011111100101100111: color_data = 12'b111100001111;
20'b01011111100101101000: color_data = 12'b111100001111;
20'b01011111100101101001: color_data = 12'b111100001111;
20'b01011111100101101010: color_data = 12'b111100001111;
20'b01011111100101101011: color_data = 12'b111100001111;
20'b01011111100101101100: color_data = 12'b111100001111;
20'b01011111100101101101: color_data = 12'b111100001111;
20'b01011111100101101110: color_data = 12'b111100001111;
20'b01011111100101101111: color_data = 12'b111100001111;
20'b01011111100101110000: color_data = 12'b111100001111;
20'b01011111100101110001: color_data = 12'b111100001111;
20'b01011111100101110010: color_data = 12'b111100001111;
20'b01011111100101110011: color_data = 12'b111100001111;
20'b01011111100101110100: color_data = 12'b111100001111;
20'b01011111100110001101: color_data = 12'b111100000000;
20'b01011111100110001110: color_data = 12'b111100000000;
20'b01011111100110001111: color_data = 12'b111100000000;
20'b01011111100110010000: color_data = 12'b111100000000;
20'b01011111100110010001: color_data = 12'b111100000000;
20'b01011111100110010010: color_data = 12'b111100000000;
20'b01011111100110010011: color_data = 12'b111100000000;
20'b01011111100110010100: color_data = 12'b111100000000;
20'b01011111100110010101: color_data = 12'b111100000000;
20'b01011111100110010110: color_data = 12'b111100000000;
20'b01011111100110010111: color_data = 12'b111100000000;
20'b01011111100110011000: color_data = 12'b111100000000;
20'b01011111100110011001: color_data = 12'b111100000000;
20'b01011111100110011010: color_data = 12'b111100000000;
20'b01011111100110011011: color_data = 12'b111100000000;
20'b01011111100110011100: color_data = 12'b111100000000;
20'b01011111100110011101: color_data = 12'b111100000000;
20'b01011111100110011110: color_data = 12'b111100000000;
20'b01011111110011111010: color_data = 12'b000011111111;
20'b01011111110011111011: color_data = 12'b000011111111;
20'b01011111110011111100: color_data = 12'b000011111111;
20'b01011111110011111101: color_data = 12'b000011111111;
20'b01011111110011111110: color_data = 12'b000011111111;
20'b01011111110011111111: color_data = 12'b000011111111;
20'b01011111110100000000: color_data = 12'b000011111111;
20'b01011111110100000001: color_data = 12'b000011111111;
20'b01011111110100000010: color_data = 12'b000011111111;
20'b01011111110100000011: color_data = 12'b000011111111;
20'b01011111110100000100: color_data = 12'b000011111111;
20'b01011111110100000101: color_data = 12'b000011111111;
20'b01011111110100000110: color_data = 12'b000011111111;
20'b01011111110100000111: color_data = 12'b000011111111;
20'b01011111110100001000: color_data = 12'b000011111111;
20'b01011111110100001001: color_data = 12'b000011111111;
20'b01011111110100001010: color_data = 12'b000011111111;
20'b01011111110100001011: color_data = 12'b000011111111;
20'b01011111110100001111: color_data = 12'b000011111111;
20'b01011111110100010000: color_data = 12'b000011111111;
20'b01011111110100010001: color_data = 12'b000011111111;
20'b01011111110100010010: color_data = 12'b000011111111;
20'b01011111110100010011: color_data = 12'b000011111111;
20'b01011111110100010100: color_data = 12'b000011111111;
20'b01011111110100010101: color_data = 12'b000011111111;
20'b01011111110100010110: color_data = 12'b000011111111;
20'b01011111110100010111: color_data = 12'b000011111111;
20'b01011111110100011000: color_data = 12'b000011111111;
20'b01011111110100011001: color_data = 12'b000011111111;
20'b01011111110100011010: color_data = 12'b000011111111;
20'b01011111110100011011: color_data = 12'b000011111111;
20'b01011111110100011100: color_data = 12'b000011111111;
20'b01011111110100011101: color_data = 12'b000011111111;
20'b01011111110100011110: color_data = 12'b000011111111;
20'b01011111110100011111: color_data = 12'b000011111111;
20'b01011111110100100000: color_data = 12'b000011111111;
20'b01011111110100100100: color_data = 12'b000001101111;
20'b01011111110100100101: color_data = 12'b000001101111;
20'b01011111110100100110: color_data = 12'b000001101111;
20'b01011111110100100111: color_data = 12'b000001101111;
20'b01011111110100101000: color_data = 12'b000001101111;
20'b01011111110100101001: color_data = 12'b000001101111;
20'b01011111110100101010: color_data = 12'b000001101111;
20'b01011111110100101011: color_data = 12'b000001101111;
20'b01011111110100101100: color_data = 12'b000001101111;
20'b01011111110100101101: color_data = 12'b000001101111;
20'b01011111110100101110: color_data = 12'b000001101111;
20'b01011111110100101111: color_data = 12'b000001101111;
20'b01011111110100110000: color_data = 12'b000001101111;
20'b01011111110100110001: color_data = 12'b000001101111;
20'b01011111110100110010: color_data = 12'b000001101111;
20'b01011111110100110011: color_data = 12'b000001101111;
20'b01011111110100110100: color_data = 12'b000001101111;
20'b01011111110100110101: color_data = 12'b000001101111;
20'b01011111110100111001: color_data = 12'b000011110000;
20'b01011111110100111010: color_data = 12'b000011110000;
20'b01011111110100111011: color_data = 12'b000011110000;
20'b01011111110100111100: color_data = 12'b000011110000;
20'b01011111110100111101: color_data = 12'b000011110000;
20'b01011111110100111110: color_data = 12'b000011110000;
20'b01011111110100111111: color_data = 12'b000011110000;
20'b01011111110101000000: color_data = 12'b000011110000;
20'b01011111110101000001: color_data = 12'b000011110000;
20'b01011111110101000010: color_data = 12'b000011110000;
20'b01011111110101000011: color_data = 12'b000011110000;
20'b01011111110101000100: color_data = 12'b000011110000;
20'b01011111110101000101: color_data = 12'b000011110000;
20'b01011111110101000110: color_data = 12'b000011110000;
20'b01011111110101000111: color_data = 12'b000011110000;
20'b01011111110101001000: color_data = 12'b000011110000;
20'b01011111110101001001: color_data = 12'b000011110000;
20'b01011111110101001010: color_data = 12'b000011110000;
20'b01011111110101100011: color_data = 12'b111100001111;
20'b01011111110101100100: color_data = 12'b111100001111;
20'b01011111110101100101: color_data = 12'b111100001111;
20'b01011111110101100110: color_data = 12'b111100001111;
20'b01011111110101100111: color_data = 12'b111100001111;
20'b01011111110101101000: color_data = 12'b111100001111;
20'b01011111110101101001: color_data = 12'b111100001111;
20'b01011111110101101010: color_data = 12'b111100001111;
20'b01011111110101101011: color_data = 12'b111100001111;
20'b01011111110101101100: color_data = 12'b111100001111;
20'b01011111110101101101: color_data = 12'b111100001111;
20'b01011111110101101110: color_data = 12'b111100001111;
20'b01011111110101101111: color_data = 12'b111100001111;
20'b01011111110101110000: color_data = 12'b111100001111;
20'b01011111110101110001: color_data = 12'b111100001111;
20'b01011111110101110010: color_data = 12'b111100001111;
20'b01011111110101110011: color_data = 12'b111100001111;
20'b01011111110101110100: color_data = 12'b111100001111;
20'b01011111110110001101: color_data = 12'b111100000000;
20'b01011111110110001110: color_data = 12'b111100000000;
20'b01011111110110001111: color_data = 12'b111100000000;
20'b01011111110110010000: color_data = 12'b111100000000;
20'b01011111110110010001: color_data = 12'b111100000000;
20'b01011111110110010010: color_data = 12'b111100000000;
20'b01011111110110010011: color_data = 12'b111100000000;
20'b01011111110110010100: color_data = 12'b111100000000;
20'b01011111110110010101: color_data = 12'b111100000000;
20'b01011111110110010110: color_data = 12'b111100000000;
20'b01011111110110010111: color_data = 12'b111100000000;
20'b01011111110110011000: color_data = 12'b111100000000;
20'b01011111110110011001: color_data = 12'b111100000000;
20'b01011111110110011010: color_data = 12'b111100000000;
20'b01011111110110011011: color_data = 12'b111100000000;
20'b01011111110110011100: color_data = 12'b111100000000;
20'b01011111110110011101: color_data = 12'b111100000000;
20'b01011111110110011110: color_data = 12'b111100000000;
20'b01100000000011111010: color_data = 12'b000011111111;
20'b01100000000011111011: color_data = 12'b000011111111;
20'b01100000000011111100: color_data = 12'b000011111111;
20'b01100000000011111101: color_data = 12'b000011111111;
20'b01100000000011111110: color_data = 12'b000011111111;
20'b01100000000011111111: color_data = 12'b000011111111;
20'b01100000000100000000: color_data = 12'b000011111111;
20'b01100000000100000001: color_data = 12'b000011111111;
20'b01100000000100000010: color_data = 12'b000011111111;
20'b01100000000100000011: color_data = 12'b000011111111;
20'b01100000000100000100: color_data = 12'b000011111111;
20'b01100000000100000101: color_data = 12'b000011111111;
20'b01100000000100000110: color_data = 12'b000011111111;
20'b01100000000100000111: color_data = 12'b000011111111;
20'b01100000000100001000: color_data = 12'b000011111111;
20'b01100000000100001001: color_data = 12'b000011111111;
20'b01100000000100001010: color_data = 12'b000011111111;
20'b01100000000100001011: color_data = 12'b000011111111;
20'b01100000000100001111: color_data = 12'b000011111111;
20'b01100000000100010000: color_data = 12'b000011111111;
20'b01100000000100010001: color_data = 12'b000011111111;
20'b01100000000100010010: color_data = 12'b000011111111;
20'b01100000000100010011: color_data = 12'b000011111111;
20'b01100000000100010100: color_data = 12'b000011111111;
20'b01100000000100010101: color_data = 12'b000011111111;
20'b01100000000100010110: color_data = 12'b000011111111;
20'b01100000000100010111: color_data = 12'b000011111111;
20'b01100000000100011000: color_data = 12'b000011111111;
20'b01100000000100011001: color_data = 12'b000011111111;
20'b01100000000100011010: color_data = 12'b000011111111;
20'b01100000000100011011: color_data = 12'b000011111111;
20'b01100000000100011100: color_data = 12'b000011111111;
20'b01100000000100011101: color_data = 12'b000011111111;
20'b01100000000100011110: color_data = 12'b000011111111;
20'b01100000000100011111: color_data = 12'b000011111111;
20'b01100000000100100000: color_data = 12'b000011111111;
20'b01100000000100100100: color_data = 12'b000001101111;
20'b01100000000100100101: color_data = 12'b000001101111;
20'b01100000000100100110: color_data = 12'b000001101111;
20'b01100000000100100111: color_data = 12'b000001101111;
20'b01100000000100101000: color_data = 12'b000001101111;
20'b01100000000100101001: color_data = 12'b000001101111;
20'b01100000000100101010: color_data = 12'b000001101111;
20'b01100000000100101011: color_data = 12'b000001101111;
20'b01100000000100101100: color_data = 12'b000001101111;
20'b01100000000100101101: color_data = 12'b000001101111;
20'b01100000000100101110: color_data = 12'b000001101111;
20'b01100000000100101111: color_data = 12'b000001101111;
20'b01100000000100110000: color_data = 12'b000001101111;
20'b01100000000100110001: color_data = 12'b000001101111;
20'b01100000000100110010: color_data = 12'b000001101111;
20'b01100000000100110011: color_data = 12'b000001101111;
20'b01100000000100110100: color_data = 12'b000001101111;
20'b01100000000100110101: color_data = 12'b000001101111;
20'b01100000000100111001: color_data = 12'b000011110000;
20'b01100000000100111010: color_data = 12'b000011110000;
20'b01100000000100111011: color_data = 12'b000011110000;
20'b01100000000100111100: color_data = 12'b000011110000;
20'b01100000000100111101: color_data = 12'b000011110000;
20'b01100000000100111110: color_data = 12'b000011110000;
20'b01100000000100111111: color_data = 12'b000011110000;
20'b01100000000101000000: color_data = 12'b000011110000;
20'b01100000000101000001: color_data = 12'b000011110000;
20'b01100000000101000010: color_data = 12'b000011110000;
20'b01100000000101000011: color_data = 12'b000011110000;
20'b01100000000101000100: color_data = 12'b000011110000;
20'b01100000000101000101: color_data = 12'b000011110000;
20'b01100000000101000110: color_data = 12'b000011110000;
20'b01100000000101000111: color_data = 12'b000011110000;
20'b01100000000101001000: color_data = 12'b000011110000;
20'b01100000000101001001: color_data = 12'b000011110000;
20'b01100000000101001010: color_data = 12'b000011110000;
20'b01100000000101100011: color_data = 12'b111100001111;
20'b01100000000101100100: color_data = 12'b111100001111;
20'b01100000000101100101: color_data = 12'b111100001111;
20'b01100000000101100110: color_data = 12'b111100001111;
20'b01100000000101100111: color_data = 12'b111100001111;
20'b01100000000101101000: color_data = 12'b111100001111;
20'b01100000000101101001: color_data = 12'b111100001111;
20'b01100000000101101010: color_data = 12'b111100001111;
20'b01100000000101101011: color_data = 12'b111100001111;
20'b01100000000101101100: color_data = 12'b111100001111;
20'b01100000000101101101: color_data = 12'b111100001111;
20'b01100000000101101110: color_data = 12'b111100001111;
20'b01100000000101101111: color_data = 12'b111100001111;
20'b01100000000101110000: color_data = 12'b111100001111;
20'b01100000000101110001: color_data = 12'b111100001111;
20'b01100000000101110010: color_data = 12'b111100001111;
20'b01100000000101110011: color_data = 12'b111100001111;
20'b01100000000101110100: color_data = 12'b111100001111;
20'b01100000000110001101: color_data = 12'b111100000000;
20'b01100000000110001110: color_data = 12'b111100000000;
20'b01100000000110001111: color_data = 12'b111100000000;
20'b01100000000110010000: color_data = 12'b111100000000;
20'b01100000000110010001: color_data = 12'b111100000000;
20'b01100000000110010010: color_data = 12'b111100000000;
20'b01100000000110010011: color_data = 12'b111100000000;
20'b01100000000110010100: color_data = 12'b111100000000;
20'b01100000000110010101: color_data = 12'b111100000000;
20'b01100000000110010110: color_data = 12'b111100000000;
20'b01100000000110010111: color_data = 12'b111100000000;
20'b01100000000110011000: color_data = 12'b111100000000;
20'b01100000000110011001: color_data = 12'b111100000000;
20'b01100000000110011010: color_data = 12'b111100000000;
20'b01100000000110011011: color_data = 12'b111100000000;
20'b01100000000110011100: color_data = 12'b111100000000;
20'b01100000000110011101: color_data = 12'b111100000000;
20'b01100000000110011110: color_data = 12'b111100000000;
20'b01100000010011111010: color_data = 12'b000011111111;
20'b01100000010011111011: color_data = 12'b000011111111;
20'b01100000010011111100: color_data = 12'b000011111111;
20'b01100000010011111101: color_data = 12'b000011111111;
20'b01100000010011111110: color_data = 12'b000011111111;
20'b01100000010011111111: color_data = 12'b000011111111;
20'b01100000010100000000: color_data = 12'b000011111111;
20'b01100000010100000001: color_data = 12'b000011111111;
20'b01100000010100000010: color_data = 12'b000011111111;
20'b01100000010100000011: color_data = 12'b000011111111;
20'b01100000010100000100: color_data = 12'b000011111111;
20'b01100000010100000101: color_data = 12'b000011111111;
20'b01100000010100000110: color_data = 12'b000011111111;
20'b01100000010100000111: color_data = 12'b000011111111;
20'b01100000010100001000: color_data = 12'b000011111111;
20'b01100000010100001001: color_data = 12'b000011111111;
20'b01100000010100001010: color_data = 12'b000011111111;
20'b01100000010100001011: color_data = 12'b000011111111;
20'b01100000010100001111: color_data = 12'b000011111111;
20'b01100000010100010000: color_data = 12'b000011111111;
20'b01100000010100010001: color_data = 12'b000011111111;
20'b01100000010100010010: color_data = 12'b000011111111;
20'b01100000010100010011: color_data = 12'b000011111111;
20'b01100000010100010100: color_data = 12'b000011111111;
20'b01100000010100010101: color_data = 12'b000011111111;
20'b01100000010100010110: color_data = 12'b000011111111;
20'b01100000010100010111: color_data = 12'b000011111111;
20'b01100000010100011000: color_data = 12'b000011111111;
20'b01100000010100011001: color_data = 12'b000011111111;
20'b01100000010100011010: color_data = 12'b000011111111;
20'b01100000010100011011: color_data = 12'b000011111111;
20'b01100000010100011100: color_data = 12'b000011111111;
20'b01100000010100011101: color_data = 12'b000011111111;
20'b01100000010100011110: color_data = 12'b000011111111;
20'b01100000010100011111: color_data = 12'b000011111111;
20'b01100000010100100000: color_data = 12'b000011111111;
20'b01100000010100100100: color_data = 12'b000001101111;
20'b01100000010100100101: color_data = 12'b000001101111;
20'b01100000010100100110: color_data = 12'b000001101111;
20'b01100000010100100111: color_data = 12'b000001101111;
20'b01100000010100101000: color_data = 12'b000001101111;
20'b01100000010100101001: color_data = 12'b000001101111;
20'b01100000010100101010: color_data = 12'b000001101111;
20'b01100000010100101011: color_data = 12'b000001101111;
20'b01100000010100101100: color_data = 12'b000001101111;
20'b01100000010100101101: color_data = 12'b000001101111;
20'b01100000010100101110: color_data = 12'b000001101111;
20'b01100000010100101111: color_data = 12'b000001101111;
20'b01100000010100110000: color_data = 12'b000001101111;
20'b01100000010100110001: color_data = 12'b000001101111;
20'b01100000010100110010: color_data = 12'b000001101111;
20'b01100000010100110011: color_data = 12'b000001101111;
20'b01100000010100110100: color_data = 12'b000001101111;
20'b01100000010100110101: color_data = 12'b000001101111;
20'b01100000010100111001: color_data = 12'b000011110000;
20'b01100000010100111010: color_data = 12'b000011110000;
20'b01100000010100111011: color_data = 12'b000011110000;
20'b01100000010100111100: color_data = 12'b000011110000;
20'b01100000010100111101: color_data = 12'b000011110000;
20'b01100000010100111110: color_data = 12'b000011110000;
20'b01100000010100111111: color_data = 12'b000011110000;
20'b01100000010101000000: color_data = 12'b000011110000;
20'b01100000010101000001: color_data = 12'b000011110000;
20'b01100000010101000010: color_data = 12'b000011110000;
20'b01100000010101000011: color_data = 12'b000011110000;
20'b01100000010101000100: color_data = 12'b000011110000;
20'b01100000010101000101: color_data = 12'b000011110000;
20'b01100000010101000110: color_data = 12'b000011110000;
20'b01100000010101000111: color_data = 12'b000011110000;
20'b01100000010101001000: color_data = 12'b000011110000;
20'b01100000010101001001: color_data = 12'b000011110000;
20'b01100000010101001010: color_data = 12'b000011110000;
20'b01100000010101100011: color_data = 12'b111100001111;
20'b01100000010101100100: color_data = 12'b111100001111;
20'b01100000010101100101: color_data = 12'b111100001111;
20'b01100000010101100110: color_data = 12'b111100001111;
20'b01100000010101100111: color_data = 12'b111100001111;
20'b01100000010101101000: color_data = 12'b111100001111;
20'b01100000010101101001: color_data = 12'b111100001111;
20'b01100000010101101010: color_data = 12'b111100001111;
20'b01100000010101101011: color_data = 12'b111100001111;
20'b01100000010101101100: color_data = 12'b111100001111;
20'b01100000010101101101: color_data = 12'b111100001111;
20'b01100000010101101110: color_data = 12'b111100001111;
20'b01100000010101101111: color_data = 12'b111100001111;
20'b01100000010101110000: color_data = 12'b111100001111;
20'b01100000010101110001: color_data = 12'b111100001111;
20'b01100000010101110010: color_data = 12'b111100001111;
20'b01100000010101110011: color_data = 12'b111100001111;
20'b01100000010101110100: color_data = 12'b111100001111;
20'b01100000010110001101: color_data = 12'b111100000000;
20'b01100000010110001110: color_data = 12'b111100000000;
20'b01100000010110001111: color_data = 12'b111100000000;
20'b01100000010110010000: color_data = 12'b111100000000;
20'b01100000010110010001: color_data = 12'b111100000000;
20'b01100000010110010010: color_data = 12'b111100000000;
20'b01100000010110010011: color_data = 12'b111100000000;
20'b01100000010110010100: color_data = 12'b111100000000;
20'b01100000010110010101: color_data = 12'b111100000000;
20'b01100000010110010110: color_data = 12'b111100000000;
20'b01100000010110010111: color_data = 12'b111100000000;
20'b01100000010110011000: color_data = 12'b111100000000;
20'b01100000010110011001: color_data = 12'b111100000000;
20'b01100000010110011010: color_data = 12'b111100000000;
20'b01100000010110011011: color_data = 12'b111100000000;
20'b01100000010110011100: color_data = 12'b111100000000;
20'b01100000010110011101: color_data = 12'b111100000000;
20'b01100000010110011110: color_data = 12'b111100000000;
20'b01100000100011111010: color_data = 12'b000011111111;
20'b01100000100011111011: color_data = 12'b000011111111;
20'b01100000100011111100: color_data = 12'b000011111111;
20'b01100000100011111101: color_data = 12'b000011111111;
20'b01100000100011111110: color_data = 12'b000011111111;
20'b01100000100011111111: color_data = 12'b000011111111;
20'b01100000100100000000: color_data = 12'b000011111111;
20'b01100000100100000001: color_data = 12'b000011111111;
20'b01100000100100000010: color_data = 12'b000011111111;
20'b01100000100100000011: color_data = 12'b000011111111;
20'b01100000100100000100: color_data = 12'b000011111111;
20'b01100000100100000101: color_data = 12'b000011111111;
20'b01100000100100000110: color_data = 12'b000011111111;
20'b01100000100100000111: color_data = 12'b000011111111;
20'b01100000100100001000: color_data = 12'b000011111111;
20'b01100000100100001001: color_data = 12'b000011111111;
20'b01100000100100001010: color_data = 12'b000011111111;
20'b01100000100100001011: color_data = 12'b000011111111;
20'b01100000100100001111: color_data = 12'b000011111111;
20'b01100000100100010000: color_data = 12'b000011111111;
20'b01100000100100010001: color_data = 12'b000011111111;
20'b01100000100100010010: color_data = 12'b000011111111;
20'b01100000100100010011: color_data = 12'b000011111111;
20'b01100000100100010100: color_data = 12'b000011111111;
20'b01100000100100010101: color_data = 12'b000011111111;
20'b01100000100100010110: color_data = 12'b000011111111;
20'b01100000100100010111: color_data = 12'b000011111111;
20'b01100000100100011000: color_data = 12'b000011111111;
20'b01100000100100011001: color_data = 12'b000011111111;
20'b01100000100100011010: color_data = 12'b000011111111;
20'b01100000100100011011: color_data = 12'b000011111111;
20'b01100000100100011100: color_data = 12'b000011111111;
20'b01100000100100011101: color_data = 12'b000011111111;
20'b01100000100100011110: color_data = 12'b000011111111;
20'b01100000100100011111: color_data = 12'b000011111111;
20'b01100000100100100000: color_data = 12'b000011111111;
20'b01100000100100100100: color_data = 12'b000001101111;
20'b01100000100100100101: color_data = 12'b000001101111;
20'b01100000100100100110: color_data = 12'b000001101111;
20'b01100000100100100111: color_data = 12'b000001101111;
20'b01100000100100101000: color_data = 12'b000001101111;
20'b01100000100100101001: color_data = 12'b000001101111;
20'b01100000100100101010: color_data = 12'b000001101111;
20'b01100000100100101011: color_data = 12'b000001101111;
20'b01100000100100101100: color_data = 12'b000001101111;
20'b01100000100100101101: color_data = 12'b000001101111;
20'b01100000100100101110: color_data = 12'b000001101111;
20'b01100000100100101111: color_data = 12'b000001101111;
20'b01100000100100110000: color_data = 12'b000001101111;
20'b01100000100100110001: color_data = 12'b000001101111;
20'b01100000100100110010: color_data = 12'b000001101111;
20'b01100000100100110011: color_data = 12'b000001101111;
20'b01100000100100110100: color_data = 12'b000001101111;
20'b01100000100100110101: color_data = 12'b000001101111;
20'b01100000100100111001: color_data = 12'b000011110000;
20'b01100000100100111010: color_data = 12'b000011110000;
20'b01100000100100111011: color_data = 12'b000011110000;
20'b01100000100100111100: color_data = 12'b000011110000;
20'b01100000100100111101: color_data = 12'b000011110000;
20'b01100000100100111110: color_data = 12'b000011110000;
20'b01100000100100111111: color_data = 12'b000011110000;
20'b01100000100101000000: color_data = 12'b000011110000;
20'b01100000100101000001: color_data = 12'b000011110000;
20'b01100000100101000010: color_data = 12'b000011110000;
20'b01100000100101000011: color_data = 12'b000011110000;
20'b01100000100101000100: color_data = 12'b000011110000;
20'b01100000100101000101: color_data = 12'b000011110000;
20'b01100000100101000110: color_data = 12'b000011110000;
20'b01100000100101000111: color_data = 12'b000011110000;
20'b01100000100101001000: color_data = 12'b000011110000;
20'b01100000100101001001: color_data = 12'b000011110000;
20'b01100000100101001010: color_data = 12'b000011110000;
20'b01100000100101100011: color_data = 12'b111100001111;
20'b01100000100101100100: color_data = 12'b111100001111;
20'b01100000100101100101: color_data = 12'b111100001111;
20'b01100000100101100110: color_data = 12'b111100001111;
20'b01100000100101100111: color_data = 12'b111100001111;
20'b01100000100101101000: color_data = 12'b111100001111;
20'b01100000100101101001: color_data = 12'b111100001111;
20'b01100000100101101010: color_data = 12'b111100001111;
20'b01100000100101101011: color_data = 12'b111100001111;
20'b01100000100101101100: color_data = 12'b111100001111;
20'b01100000100101101101: color_data = 12'b111100001111;
20'b01100000100101101110: color_data = 12'b111100001111;
20'b01100000100101101111: color_data = 12'b111100001111;
20'b01100000100101110000: color_data = 12'b111100001111;
20'b01100000100101110001: color_data = 12'b111100001111;
20'b01100000100101110010: color_data = 12'b111100001111;
20'b01100000100101110011: color_data = 12'b111100001111;
20'b01100000100101110100: color_data = 12'b111100001111;
20'b01100000100110001101: color_data = 12'b111100000000;
20'b01100000100110001110: color_data = 12'b111100000000;
20'b01100000100110001111: color_data = 12'b111100000000;
20'b01100000100110010000: color_data = 12'b111100000000;
20'b01100000100110010001: color_data = 12'b111100000000;
20'b01100000100110010010: color_data = 12'b111100000000;
20'b01100000100110010011: color_data = 12'b111100000000;
20'b01100000100110010100: color_data = 12'b111100000000;
20'b01100000100110010101: color_data = 12'b111100000000;
20'b01100000100110010110: color_data = 12'b111100000000;
20'b01100000100110010111: color_data = 12'b111100000000;
20'b01100000100110011000: color_data = 12'b111100000000;
20'b01100000100110011001: color_data = 12'b111100000000;
20'b01100000100110011010: color_data = 12'b111100000000;
20'b01100000100110011011: color_data = 12'b111100000000;
20'b01100000100110011100: color_data = 12'b111100000000;
20'b01100000100110011101: color_data = 12'b111100000000;
20'b01100000100110011110: color_data = 12'b111100000000;
20'b01100000110011111010: color_data = 12'b000011111111;
20'b01100000110011111011: color_data = 12'b000011111111;
20'b01100000110011111100: color_data = 12'b000011111111;
20'b01100000110011111101: color_data = 12'b000011111111;
20'b01100000110011111110: color_data = 12'b000011111111;
20'b01100000110011111111: color_data = 12'b000011111111;
20'b01100000110100000000: color_data = 12'b000011111111;
20'b01100000110100000001: color_data = 12'b000011111111;
20'b01100000110100000010: color_data = 12'b000011111111;
20'b01100000110100000011: color_data = 12'b000011111111;
20'b01100000110100000100: color_data = 12'b000011111111;
20'b01100000110100000101: color_data = 12'b000011111111;
20'b01100000110100000110: color_data = 12'b000011111111;
20'b01100000110100000111: color_data = 12'b000011111111;
20'b01100000110100001000: color_data = 12'b000011111111;
20'b01100000110100001001: color_data = 12'b000011111111;
20'b01100000110100001010: color_data = 12'b000011111111;
20'b01100000110100001011: color_data = 12'b000011111111;
20'b01100000110100001111: color_data = 12'b000011111111;
20'b01100000110100010000: color_data = 12'b000011111111;
20'b01100000110100010001: color_data = 12'b000011111111;
20'b01100000110100010010: color_data = 12'b000011111111;
20'b01100000110100010011: color_data = 12'b000011111111;
20'b01100000110100010100: color_data = 12'b000011111111;
20'b01100000110100010101: color_data = 12'b000011111111;
20'b01100000110100010110: color_data = 12'b000011111111;
20'b01100000110100010111: color_data = 12'b000011111111;
20'b01100000110100011000: color_data = 12'b000011111111;
20'b01100000110100011001: color_data = 12'b000011111111;
20'b01100000110100011010: color_data = 12'b000011111111;
20'b01100000110100011011: color_data = 12'b000011111111;
20'b01100000110100011100: color_data = 12'b000011111111;
20'b01100000110100011101: color_data = 12'b000011111111;
20'b01100000110100011110: color_data = 12'b000011111111;
20'b01100000110100011111: color_data = 12'b000011111111;
20'b01100000110100100000: color_data = 12'b000011111111;
20'b01100000110100100100: color_data = 12'b000001101111;
20'b01100000110100100101: color_data = 12'b000001101111;
20'b01100000110100100110: color_data = 12'b000001101111;
20'b01100000110100100111: color_data = 12'b000001101111;
20'b01100000110100101000: color_data = 12'b000001101111;
20'b01100000110100101001: color_data = 12'b000001101111;
20'b01100000110100101010: color_data = 12'b000001101111;
20'b01100000110100101011: color_data = 12'b000001101111;
20'b01100000110100101100: color_data = 12'b000001101111;
20'b01100000110100101101: color_data = 12'b000001101111;
20'b01100000110100101110: color_data = 12'b000001101111;
20'b01100000110100101111: color_data = 12'b000001101111;
20'b01100000110100110000: color_data = 12'b000001101111;
20'b01100000110100110001: color_data = 12'b000001101111;
20'b01100000110100110010: color_data = 12'b000001101111;
20'b01100000110100110011: color_data = 12'b000001101111;
20'b01100000110100110100: color_data = 12'b000001101111;
20'b01100000110100110101: color_data = 12'b000001101111;
20'b01100000110100111001: color_data = 12'b000011110000;
20'b01100000110100111010: color_data = 12'b000011110000;
20'b01100000110100111011: color_data = 12'b000011110000;
20'b01100000110100111100: color_data = 12'b000011110000;
20'b01100000110100111101: color_data = 12'b000011110000;
20'b01100000110100111110: color_data = 12'b000011110000;
20'b01100000110100111111: color_data = 12'b000011110000;
20'b01100000110101000000: color_data = 12'b000011110000;
20'b01100000110101000001: color_data = 12'b000011110000;
20'b01100000110101000010: color_data = 12'b000011110000;
20'b01100000110101000011: color_data = 12'b000011110000;
20'b01100000110101000100: color_data = 12'b000011110000;
20'b01100000110101000101: color_data = 12'b000011110000;
20'b01100000110101000110: color_data = 12'b000011110000;
20'b01100000110101000111: color_data = 12'b000011110000;
20'b01100000110101001000: color_data = 12'b000011110000;
20'b01100000110101001001: color_data = 12'b000011110000;
20'b01100000110101001010: color_data = 12'b000011110000;
20'b01100000110101100011: color_data = 12'b111100001111;
20'b01100000110101100100: color_data = 12'b111100001111;
20'b01100000110101100101: color_data = 12'b111100001111;
20'b01100000110101100110: color_data = 12'b111100001111;
20'b01100000110101100111: color_data = 12'b111100001111;
20'b01100000110101101000: color_data = 12'b111100001111;
20'b01100000110101101001: color_data = 12'b111100001111;
20'b01100000110101101010: color_data = 12'b111100001111;
20'b01100000110101101011: color_data = 12'b111100001111;
20'b01100000110101101100: color_data = 12'b111100001111;
20'b01100000110101101101: color_data = 12'b111100001111;
20'b01100000110101101110: color_data = 12'b111100001111;
20'b01100000110101101111: color_data = 12'b111100001111;
20'b01100000110101110000: color_data = 12'b111100001111;
20'b01100000110101110001: color_data = 12'b111100001111;
20'b01100000110101110010: color_data = 12'b111100001111;
20'b01100000110101110011: color_data = 12'b111100001111;
20'b01100000110101110100: color_data = 12'b111100001111;
20'b01100000110110001101: color_data = 12'b111100000000;
20'b01100000110110001110: color_data = 12'b111100000000;
20'b01100000110110001111: color_data = 12'b111100000000;
20'b01100000110110010000: color_data = 12'b111100000000;
20'b01100000110110010001: color_data = 12'b111100000000;
20'b01100000110110010010: color_data = 12'b111100000000;
20'b01100000110110010011: color_data = 12'b111100000000;
20'b01100000110110010100: color_data = 12'b111100000000;
20'b01100000110110010101: color_data = 12'b111100000000;
20'b01100000110110010110: color_data = 12'b111100000000;
20'b01100000110110010111: color_data = 12'b111100000000;
20'b01100000110110011000: color_data = 12'b111100000000;
20'b01100000110110011001: color_data = 12'b111100000000;
20'b01100000110110011010: color_data = 12'b111100000000;
20'b01100000110110011011: color_data = 12'b111100000000;
20'b01100000110110011100: color_data = 12'b111100000000;
20'b01100000110110011101: color_data = 12'b111100000000;
20'b01100000110110011110: color_data = 12'b111100000000;
20'b01100001000011111010: color_data = 12'b000011111111;
20'b01100001000011111011: color_data = 12'b000011111111;
20'b01100001000011111100: color_data = 12'b000011111111;
20'b01100001000011111101: color_data = 12'b000011111111;
20'b01100001000011111110: color_data = 12'b000011111111;
20'b01100001000011111111: color_data = 12'b000011111111;
20'b01100001000100000000: color_data = 12'b000011111111;
20'b01100001000100000001: color_data = 12'b000011111111;
20'b01100001000100000010: color_data = 12'b000011111111;
20'b01100001000100000011: color_data = 12'b000011111111;
20'b01100001000100000100: color_data = 12'b000011111111;
20'b01100001000100000101: color_data = 12'b000011111111;
20'b01100001000100000110: color_data = 12'b000011111111;
20'b01100001000100000111: color_data = 12'b000011111111;
20'b01100001000100001000: color_data = 12'b000011111111;
20'b01100001000100001001: color_data = 12'b000011111111;
20'b01100001000100001010: color_data = 12'b000011111111;
20'b01100001000100001011: color_data = 12'b000011111111;
20'b01100001000100001111: color_data = 12'b000011111111;
20'b01100001000100010000: color_data = 12'b000011111111;
20'b01100001000100010001: color_data = 12'b000011111111;
20'b01100001000100010010: color_data = 12'b000011111111;
20'b01100001000100010011: color_data = 12'b000011111111;
20'b01100001000100010100: color_data = 12'b000011111111;
20'b01100001000100010101: color_data = 12'b000011111111;
20'b01100001000100010110: color_data = 12'b000011111111;
20'b01100001000100010111: color_data = 12'b000011111111;
20'b01100001000100011000: color_data = 12'b000011111111;
20'b01100001000100011001: color_data = 12'b000011111111;
20'b01100001000100011010: color_data = 12'b000011111111;
20'b01100001000100011011: color_data = 12'b000011111111;
20'b01100001000100011100: color_data = 12'b000011111111;
20'b01100001000100011101: color_data = 12'b000011111111;
20'b01100001000100011110: color_data = 12'b000011111111;
20'b01100001000100011111: color_data = 12'b000011111111;
20'b01100001000100100000: color_data = 12'b000011111111;
20'b01100001000100100100: color_data = 12'b000001101111;
20'b01100001000100100101: color_data = 12'b000001101111;
20'b01100001000100100110: color_data = 12'b000001101111;
20'b01100001000100100111: color_data = 12'b000001101111;
20'b01100001000100101000: color_data = 12'b000001101111;
20'b01100001000100101001: color_data = 12'b000001101111;
20'b01100001000100101010: color_data = 12'b000001101111;
20'b01100001000100101011: color_data = 12'b000001101111;
20'b01100001000100101100: color_data = 12'b000001101111;
20'b01100001000100101101: color_data = 12'b000001101111;
20'b01100001000100101110: color_data = 12'b000001101111;
20'b01100001000100101111: color_data = 12'b000001101111;
20'b01100001000100110000: color_data = 12'b000001101111;
20'b01100001000100110001: color_data = 12'b000001101111;
20'b01100001000100110010: color_data = 12'b000001101111;
20'b01100001000100110011: color_data = 12'b000001101111;
20'b01100001000100110100: color_data = 12'b000001101111;
20'b01100001000100110101: color_data = 12'b000001101111;
20'b01100001000100111001: color_data = 12'b000011110000;
20'b01100001000100111010: color_data = 12'b000011110000;
20'b01100001000100111011: color_data = 12'b000011110000;
20'b01100001000100111100: color_data = 12'b000011110000;
20'b01100001000100111101: color_data = 12'b000011110000;
20'b01100001000100111110: color_data = 12'b000011110000;
20'b01100001000100111111: color_data = 12'b000011110000;
20'b01100001000101000000: color_data = 12'b000011110000;
20'b01100001000101000001: color_data = 12'b000011110000;
20'b01100001000101000010: color_data = 12'b000011110000;
20'b01100001000101000011: color_data = 12'b000011110000;
20'b01100001000101000100: color_data = 12'b000011110000;
20'b01100001000101000101: color_data = 12'b000011110000;
20'b01100001000101000110: color_data = 12'b000011110000;
20'b01100001000101000111: color_data = 12'b000011110000;
20'b01100001000101001000: color_data = 12'b000011110000;
20'b01100001000101001001: color_data = 12'b000011110000;
20'b01100001000101001010: color_data = 12'b000011110000;
20'b01100001000101100011: color_data = 12'b111100001111;
20'b01100001000101100100: color_data = 12'b111100001111;
20'b01100001000101100101: color_data = 12'b111100001111;
20'b01100001000101100110: color_data = 12'b111100001111;
20'b01100001000101100111: color_data = 12'b111100001111;
20'b01100001000101101000: color_data = 12'b111100001111;
20'b01100001000101101001: color_data = 12'b111100001111;
20'b01100001000101101010: color_data = 12'b111100001111;
20'b01100001000101101011: color_data = 12'b111100001111;
20'b01100001000101101100: color_data = 12'b111100001111;
20'b01100001000101101101: color_data = 12'b111100001111;
20'b01100001000101101110: color_data = 12'b111100001111;
20'b01100001000101101111: color_data = 12'b111100001111;
20'b01100001000101110000: color_data = 12'b111100001111;
20'b01100001000101110001: color_data = 12'b111100001111;
20'b01100001000101110010: color_data = 12'b111100001111;
20'b01100001000101110011: color_data = 12'b111100001111;
20'b01100001000101110100: color_data = 12'b111100001111;
20'b01100001000110001101: color_data = 12'b111100000000;
20'b01100001000110001110: color_data = 12'b111100000000;
20'b01100001000110001111: color_data = 12'b111100000000;
20'b01100001000110010000: color_data = 12'b111100000000;
20'b01100001000110010001: color_data = 12'b111100000000;
20'b01100001000110010010: color_data = 12'b111100000000;
20'b01100001000110010011: color_data = 12'b111100000000;
20'b01100001000110010100: color_data = 12'b111100000000;
20'b01100001000110010101: color_data = 12'b111100000000;
20'b01100001000110010110: color_data = 12'b111100000000;
20'b01100001000110010111: color_data = 12'b111100000000;
20'b01100001000110011000: color_data = 12'b111100000000;
20'b01100001000110011001: color_data = 12'b111100000000;
20'b01100001000110011010: color_data = 12'b111100000000;
20'b01100001000110011011: color_data = 12'b111100000000;
20'b01100001000110011100: color_data = 12'b111100000000;
20'b01100001000110011101: color_data = 12'b111100000000;
20'b01100001000110011110: color_data = 12'b111100000000;
20'b01100001010011111010: color_data = 12'b000011111111;
20'b01100001010011111011: color_data = 12'b000011111111;
20'b01100001010011111100: color_data = 12'b000011111111;
20'b01100001010011111101: color_data = 12'b000011111111;
20'b01100001010011111110: color_data = 12'b000011111111;
20'b01100001010011111111: color_data = 12'b000011111111;
20'b01100001010100000000: color_data = 12'b000011111111;
20'b01100001010100000001: color_data = 12'b000011111111;
20'b01100001010100000010: color_data = 12'b000011111111;
20'b01100001010100000011: color_data = 12'b000011111111;
20'b01100001010100000100: color_data = 12'b000011111111;
20'b01100001010100000101: color_data = 12'b000011111111;
20'b01100001010100000110: color_data = 12'b000011111111;
20'b01100001010100000111: color_data = 12'b000011111111;
20'b01100001010100001000: color_data = 12'b000011111111;
20'b01100001010100001001: color_data = 12'b000011111111;
20'b01100001010100001010: color_data = 12'b000011111111;
20'b01100001010100001011: color_data = 12'b000011111111;
20'b01100001010100001111: color_data = 12'b000011111111;
20'b01100001010100010000: color_data = 12'b000011111111;
20'b01100001010100010001: color_data = 12'b000011111111;
20'b01100001010100010010: color_data = 12'b000011111111;
20'b01100001010100010011: color_data = 12'b000011111111;
20'b01100001010100010100: color_data = 12'b000011111111;
20'b01100001010100010101: color_data = 12'b000011111111;
20'b01100001010100010110: color_data = 12'b000011111111;
20'b01100001010100010111: color_data = 12'b000011111111;
20'b01100001010100011000: color_data = 12'b000011111111;
20'b01100001010100011001: color_data = 12'b000011111111;
20'b01100001010100011010: color_data = 12'b000011111111;
20'b01100001010100011011: color_data = 12'b000011111111;
20'b01100001010100011100: color_data = 12'b000011111111;
20'b01100001010100011101: color_data = 12'b000011111111;
20'b01100001010100011110: color_data = 12'b000011111111;
20'b01100001010100011111: color_data = 12'b000011111111;
20'b01100001010100100000: color_data = 12'b000011111111;
20'b01100001010100100100: color_data = 12'b000001101111;
20'b01100001010100100101: color_data = 12'b000001101111;
20'b01100001010100100110: color_data = 12'b000001101111;
20'b01100001010100100111: color_data = 12'b000001101111;
20'b01100001010100101000: color_data = 12'b000001101111;
20'b01100001010100101001: color_data = 12'b000001101111;
20'b01100001010100101010: color_data = 12'b000001101111;
20'b01100001010100101011: color_data = 12'b000001101111;
20'b01100001010100101100: color_data = 12'b000001101111;
20'b01100001010100101101: color_data = 12'b000001101111;
20'b01100001010100101110: color_data = 12'b000001101111;
20'b01100001010100101111: color_data = 12'b000001101111;
20'b01100001010100110000: color_data = 12'b000001101111;
20'b01100001010100110001: color_data = 12'b000001101111;
20'b01100001010100110010: color_data = 12'b000001101111;
20'b01100001010100110011: color_data = 12'b000001101111;
20'b01100001010100110100: color_data = 12'b000001101111;
20'b01100001010100110101: color_data = 12'b000001101111;
20'b01100001010100111001: color_data = 12'b000011110000;
20'b01100001010100111010: color_data = 12'b000011110000;
20'b01100001010100111011: color_data = 12'b000011110000;
20'b01100001010100111100: color_data = 12'b000011110000;
20'b01100001010100111101: color_data = 12'b000011110000;
20'b01100001010100111110: color_data = 12'b000011110000;
20'b01100001010100111111: color_data = 12'b000011110000;
20'b01100001010101000000: color_data = 12'b000011110000;
20'b01100001010101000001: color_data = 12'b000011110000;
20'b01100001010101000010: color_data = 12'b000011110000;
20'b01100001010101000011: color_data = 12'b000011110000;
20'b01100001010101000100: color_data = 12'b000011110000;
20'b01100001010101000101: color_data = 12'b000011110000;
20'b01100001010101000110: color_data = 12'b000011110000;
20'b01100001010101000111: color_data = 12'b000011110000;
20'b01100001010101001000: color_data = 12'b000011110000;
20'b01100001010101001001: color_data = 12'b000011110000;
20'b01100001010101001010: color_data = 12'b000011110000;
20'b01100001010101100011: color_data = 12'b111100001111;
20'b01100001010101100100: color_data = 12'b111100001111;
20'b01100001010101100101: color_data = 12'b111100001111;
20'b01100001010101100110: color_data = 12'b111100001111;
20'b01100001010101100111: color_data = 12'b111100001111;
20'b01100001010101101000: color_data = 12'b111100001111;
20'b01100001010101101001: color_data = 12'b111100001111;
20'b01100001010101101010: color_data = 12'b111100001111;
20'b01100001010101101011: color_data = 12'b111100001111;
20'b01100001010101101100: color_data = 12'b111100001111;
20'b01100001010101101101: color_data = 12'b111100001111;
20'b01100001010101101110: color_data = 12'b111100001111;
20'b01100001010101101111: color_data = 12'b111100001111;
20'b01100001010101110000: color_data = 12'b111100001111;
20'b01100001010101110001: color_data = 12'b111100001111;
20'b01100001010101110010: color_data = 12'b111100001111;
20'b01100001010101110011: color_data = 12'b111100001111;
20'b01100001010101110100: color_data = 12'b111100001111;
20'b01100001010110001101: color_data = 12'b111100000000;
20'b01100001010110001110: color_data = 12'b111100000000;
20'b01100001010110001111: color_data = 12'b111100000000;
20'b01100001010110010000: color_data = 12'b111100000000;
20'b01100001010110010001: color_data = 12'b111100000000;
20'b01100001010110010010: color_data = 12'b111100000000;
20'b01100001010110010011: color_data = 12'b111100000000;
20'b01100001010110010100: color_data = 12'b111100000000;
20'b01100001010110010101: color_data = 12'b111100000000;
20'b01100001010110010110: color_data = 12'b111100000000;
20'b01100001010110010111: color_data = 12'b111100000000;
20'b01100001010110011000: color_data = 12'b111100000000;
20'b01100001010110011001: color_data = 12'b111100000000;
20'b01100001010110011010: color_data = 12'b111100000000;
20'b01100001010110011011: color_data = 12'b111100000000;
20'b01100001010110011100: color_data = 12'b111100000000;
20'b01100001010110011101: color_data = 12'b111100000000;
20'b01100001010110011110: color_data = 12'b111100000000;
20'b01100001100011111010: color_data = 12'b000011111111;
20'b01100001100011111011: color_data = 12'b000011111111;
20'b01100001100011111100: color_data = 12'b000011111111;
20'b01100001100011111101: color_data = 12'b000011111111;
20'b01100001100011111110: color_data = 12'b000011111111;
20'b01100001100011111111: color_data = 12'b000011111111;
20'b01100001100100000000: color_data = 12'b000011111111;
20'b01100001100100000001: color_data = 12'b000011111111;
20'b01100001100100000010: color_data = 12'b000011111111;
20'b01100001100100000011: color_data = 12'b000011111111;
20'b01100001100100000100: color_data = 12'b000011111111;
20'b01100001100100000101: color_data = 12'b000011111111;
20'b01100001100100000110: color_data = 12'b000011111111;
20'b01100001100100000111: color_data = 12'b000011111111;
20'b01100001100100001000: color_data = 12'b000011111111;
20'b01100001100100001001: color_data = 12'b000011111111;
20'b01100001100100001010: color_data = 12'b000011111111;
20'b01100001100100001011: color_data = 12'b000011111111;
20'b01100001100100001111: color_data = 12'b000011111111;
20'b01100001100100010000: color_data = 12'b000011111111;
20'b01100001100100010001: color_data = 12'b000011111111;
20'b01100001100100010010: color_data = 12'b000011111111;
20'b01100001100100010011: color_data = 12'b000011111111;
20'b01100001100100010100: color_data = 12'b000011111111;
20'b01100001100100010101: color_data = 12'b000011111111;
20'b01100001100100010110: color_data = 12'b000011111111;
20'b01100001100100010111: color_data = 12'b000011111111;
20'b01100001100100011000: color_data = 12'b000011111111;
20'b01100001100100011001: color_data = 12'b000011111111;
20'b01100001100100011010: color_data = 12'b000011111111;
20'b01100001100100011011: color_data = 12'b000011111111;
20'b01100001100100011100: color_data = 12'b000011111111;
20'b01100001100100011101: color_data = 12'b000011111111;
20'b01100001100100011110: color_data = 12'b000011111111;
20'b01100001100100011111: color_data = 12'b000011111111;
20'b01100001100100100000: color_data = 12'b000011111111;
20'b01100001100100100100: color_data = 12'b000001101111;
20'b01100001100100100101: color_data = 12'b000001101111;
20'b01100001100100100110: color_data = 12'b000001101111;
20'b01100001100100100111: color_data = 12'b000001101111;
20'b01100001100100101000: color_data = 12'b000001101111;
20'b01100001100100101001: color_data = 12'b000001101111;
20'b01100001100100101010: color_data = 12'b000001101111;
20'b01100001100100101011: color_data = 12'b000001101111;
20'b01100001100100101100: color_data = 12'b000001101111;
20'b01100001100100101101: color_data = 12'b000001101111;
20'b01100001100100101110: color_data = 12'b000001101111;
20'b01100001100100101111: color_data = 12'b000001101111;
20'b01100001100100110000: color_data = 12'b000001101111;
20'b01100001100100110001: color_data = 12'b000001101111;
20'b01100001100100110010: color_data = 12'b000001101111;
20'b01100001100100110011: color_data = 12'b000001101111;
20'b01100001100100110100: color_data = 12'b000001101111;
20'b01100001100100110101: color_data = 12'b000001101111;
20'b01100001100100111001: color_data = 12'b000011110000;
20'b01100001100100111010: color_data = 12'b000011110000;
20'b01100001100100111011: color_data = 12'b000011110000;
20'b01100001100100111100: color_data = 12'b000011110000;
20'b01100001100100111101: color_data = 12'b000011110000;
20'b01100001100100111110: color_data = 12'b000011110000;
20'b01100001100100111111: color_data = 12'b000011110000;
20'b01100001100101000000: color_data = 12'b000011110000;
20'b01100001100101000001: color_data = 12'b000011110000;
20'b01100001100101000010: color_data = 12'b000011110000;
20'b01100001100101000011: color_data = 12'b000011110000;
20'b01100001100101000100: color_data = 12'b000011110000;
20'b01100001100101000101: color_data = 12'b000011110000;
20'b01100001100101000110: color_data = 12'b000011110000;
20'b01100001100101000111: color_data = 12'b000011110000;
20'b01100001100101001000: color_data = 12'b000011110000;
20'b01100001100101001001: color_data = 12'b000011110000;
20'b01100001100101001010: color_data = 12'b000011110000;
20'b01100001100101100011: color_data = 12'b111100001111;
20'b01100001100101100100: color_data = 12'b111100001111;
20'b01100001100101100101: color_data = 12'b111100001111;
20'b01100001100101100110: color_data = 12'b111100001111;
20'b01100001100101100111: color_data = 12'b111100001111;
20'b01100001100101101000: color_data = 12'b111100001111;
20'b01100001100101101001: color_data = 12'b111100001111;
20'b01100001100101101010: color_data = 12'b111100001111;
20'b01100001100101101011: color_data = 12'b111100001111;
20'b01100001100101101100: color_data = 12'b111100001111;
20'b01100001100101101101: color_data = 12'b111100001111;
20'b01100001100101101110: color_data = 12'b111100001111;
20'b01100001100101101111: color_data = 12'b111100001111;
20'b01100001100101110000: color_data = 12'b111100001111;
20'b01100001100101110001: color_data = 12'b111100001111;
20'b01100001100101110010: color_data = 12'b111100001111;
20'b01100001100101110011: color_data = 12'b111100001111;
20'b01100001100101110100: color_data = 12'b111100001111;
20'b01100001100110001101: color_data = 12'b111100000000;
20'b01100001100110001110: color_data = 12'b111100000000;
20'b01100001100110001111: color_data = 12'b111100000000;
20'b01100001100110010000: color_data = 12'b111100000000;
20'b01100001100110010001: color_data = 12'b111100000000;
20'b01100001100110010010: color_data = 12'b111100000000;
20'b01100001100110010011: color_data = 12'b111100000000;
20'b01100001100110010100: color_data = 12'b111100000000;
20'b01100001100110010101: color_data = 12'b111100000000;
20'b01100001100110010110: color_data = 12'b111100000000;
20'b01100001100110010111: color_data = 12'b111100000000;
20'b01100001100110011000: color_data = 12'b111100000000;
20'b01100001100110011001: color_data = 12'b111100000000;
20'b01100001100110011010: color_data = 12'b111100000000;
20'b01100001100110011011: color_data = 12'b111100000000;
20'b01100001100110011100: color_data = 12'b111100000000;
20'b01100001100110011101: color_data = 12'b111100000000;
20'b01100001100110011110: color_data = 12'b111100000000;
20'b01100001110011111010: color_data = 12'b000011111111;
20'b01100001110011111011: color_data = 12'b000011111111;
20'b01100001110011111100: color_data = 12'b000011111111;
20'b01100001110011111101: color_data = 12'b000011111111;
20'b01100001110011111110: color_data = 12'b000011111111;
20'b01100001110011111111: color_data = 12'b000011111111;
20'b01100001110100000000: color_data = 12'b000011111111;
20'b01100001110100000001: color_data = 12'b000011111111;
20'b01100001110100000010: color_data = 12'b000011111111;
20'b01100001110100000011: color_data = 12'b000011111111;
20'b01100001110100000100: color_data = 12'b000011111111;
20'b01100001110100000101: color_data = 12'b000011111111;
20'b01100001110100000110: color_data = 12'b000011111111;
20'b01100001110100000111: color_data = 12'b000011111111;
20'b01100001110100001000: color_data = 12'b000011111111;
20'b01100001110100001001: color_data = 12'b000011111111;
20'b01100001110100001010: color_data = 12'b000011111111;
20'b01100001110100001011: color_data = 12'b000011111111;
20'b01100001110100001111: color_data = 12'b000011111111;
20'b01100001110100010000: color_data = 12'b000011111111;
20'b01100001110100010001: color_data = 12'b000011111111;
20'b01100001110100010010: color_data = 12'b000011111111;
20'b01100001110100010011: color_data = 12'b000011111111;
20'b01100001110100010100: color_data = 12'b000011111111;
20'b01100001110100010101: color_data = 12'b000011111111;
20'b01100001110100010110: color_data = 12'b000011111111;
20'b01100001110100010111: color_data = 12'b000011111111;
20'b01100001110100011000: color_data = 12'b000011111111;
20'b01100001110100011001: color_data = 12'b000011111111;
20'b01100001110100011010: color_data = 12'b000011111111;
20'b01100001110100011011: color_data = 12'b000011111111;
20'b01100001110100011100: color_data = 12'b000011111111;
20'b01100001110100011101: color_data = 12'b000011111111;
20'b01100001110100011110: color_data = 12'b000011111111;
20'b01100001110100011111: color_data = 12'b000011111111;
20'b01100001110100100000: color_data = 12'b000011111111;
20'b01100001110100100100: color_data = 12'b000001101111;
20'b01100001110100100101: color_data = 12'b000001101111;
20'b01100001110100100110: color_data = 12'b000001101111;
20'b01100001110100100111: color_data = 12'b000001101111;
20'b01100001110100101000: color_data = 12'b000001101111;
20'b01100001110100101001: color_data = 12'b000001101111;
20'b01100001110100101010: color_data = 12'b000001101111;
20'b01100001110100101011: color_data = 12'b000001101111;
20'b01100001110100101100: color_data = 12'b000001101111;
20'b01100001110100101101: color_data = 12'b000001101111;
20'b01100001110100101110: color_data = 12'b000001101111;
20'b01100001110100101111: color_data = 12'b000001101111;
20'b01100001110100110000: color_data = 12'b000001101111;
20'b01100001110100110001: color_data = 12'b000001101111;
20'b01100001110100110010: color_data = 12'b000001101111;
20'b01100001110100110011: color_data = 12'b000001101111;
20'b01100001110100110100: color_data = 12'b000001101111;
20'b01100001110100110101: color_data = 12'b000001101111;
20'b01100001110100111001: color_data = 12'b000011110000;
20'b01100001110100111010: color_data = 12'b000011110000;
20'b01100001110100111011: color_data = 12'b000011110000;
20'b01100001110100111100: color_data = 12'b000011110000;
20'b01100001110100111101: color_data = 12'b000011110000;
20'b01100001110100111110: color_data = 12'b000011110000;
20'b01100001110100111111: color_data = 12'b000011110000;
20'b01100001110101000000: color_data = 12'b000011110000;
20'b01100001110101000001: color_data = 12'b000011110000;
20'b01100001110101000010: color_data = 12'b000011110000;
20'b01100001110101000011: color_data = 12'b000011110000;
20'b01100001110101000100: color_data = 12'b000011110000;
20'b01100001110101000101: color_data = 12'b000011110000;
20'b01100001110101000110: color_data = 12'b000011110000;
20'b01100001110101000111: color_data = 12'b000011110000;
20'b01100001110101001000: color_data = 12'b000011110000;
20'b01100001110101001001: color_data = 12'b000011110000;
20'b01100001110101001010: color_data = 12'b000011110000;
20'b01100001110101100011: color_data = 12'b111100001111;
20'b01100001110101100100: color_data = 12'b111100001111;
20'b01100001110101100101: color_data = 12'b111100001111;
20'b01100001110101100110: color_data = 12'b111100001111;
20'b01100001110101100111: color_data = 12'b111100001111;
20'b01100001110101101000: color_data = 12'b111100001111;
20'b01100001110101101001: color_data = 12'b111100001111;
20'b01100001110101101010: color_data = 12'b111100001111;
20'b01100001110101101011: color_data = 12'b111100001111;
20'b01100001110101101100: color_data = 12'b111100001111;
20'b01100001110101101101: color_data = 12'b111100001111;
20'b01100001110101101110: color_data = 12'b111100001111;
20'b01100001110101101111: color_data = 12'b111100001111;
20'b01100001110101110000: color_data = 12'b111100001111;
20'b01100001110101110001: color_data = 12'b111100001111;
20'b01100001110101110010: color_data = 12'b111100001111;
20'b01100001110101110011: color_data = 12'b111100001111;
20'b01100001110101110100: color_data = 12'b111100001111;
20'b01100001110110001101: color_data = 12'b111100000000;
20'b01100001110110001110: color_data = 12'b111100000000;
20'b01100001110110001111: color_data = 12'b111100000000;
20'b01100001110110010000: color_data = 12'b111100000000;
20'b01100001110110010001: color_data = 12'b111100000000;
20'b01100001110110010010: color_data = 12'b111100000000;
20'b01100001110110010011: color_data = 12'b111100000000;
20'b01100001110110010100: color_data = 12'b111100000000;
20'b01100001110110010101: color_data = 12'b111100000000;
20'b01100001110110010110: color_data = 12'b111100000000;
20'b01100001110110010111: color_data = 12'b111100000000;
20'b01100001110110011000: color_data = 12'b111100000000;
20'b01100001110110011001: color_data = 12'b111100000000;
20'b01100001110110011010: color_data = 12'b111100000000;
20'b01100001110110011011: color_data = 12'b111100000000;
20'b01100001110110011100: color_data = 12'b111100000000;
20'b01100001110110011101: color_data = 12'b111100000000;
20'b01100001110110011110: color_data = 12'b111100000000;
20'b01100010000011111010: color_data = 12'b000011111111;
20'b01100010000011111011: color_data = 12'b000011111111;
20'b01100010000011111100: color_data = 12'b000011111111;
20'b01100010000011111101: color_data = 12'b000011111111;
20'b01100010000011111110: color_data = 12'b000011111111;
20'b01100010000011111111: color_data = 12'b000011111111;
20'b01100010000100000000: color_data = 12'b000011111111;
20'b01100010000100000001: color_data = 12'b000011111111;
20'b01100010000100000010: color_data = 12'b000011111111;
20'b01100010000100000011: color_data = 12'b000011111111;
20'b01100010000100000100: color_data = 12'b000011111111;
20'b01100010000100000101: color_data = 12'b000011111111;
20'b01100010000100000110: color_data = 12'b000011111111;
20'b01100010000100000111: color_data = 12'b000011111111;
20'b01100010000100001000: color_data = 12'b000011111111;
20'b01100010000100001001: color_data = 12'b000011111111;
20'b01100010000100001010: color_data = 12'b000011111111;
20'b01100010000100001011: color_data = 12'b000011111111;
20'b01100010000100001111: color_data = 12'b000011111111;
20'b01100010000100010000: color_data = 12'b000011111111;
20'b01100010000100010001: color_data = 12'b000011111111;
20'b01100010000100010010: color_data = 12'b000011111111;
20'b01100010000100010011: color_data = 12'b000011111111;
20'b01100010000100010100: color_data = 12'b000011111111;
20'b01100010000100010101: color_data = 12'b000011111111;
20'b01100010000100010110: color_data = 12'b000011111111;
20'b01100010000100010111: color_data = 12'b000011111111;
20'b01100010000100011000: color_data = 12'b000011111111;
20'b01100010000100011001: color_data = 12'b000011111111;
20'b01100010000100011010: color_data = 12'b000011111111;
20'b01100010000100011011: color_data = 12'b000011111111;
20'b01100010000100011100: color_data = 12'b000011111111;
20'b01100010000100011101: color_data = 12'b000011111111;
20'b01100010000100011110: color_data = 12'b000011111111;
20'b01100010000100011111: color_data = 12'b000011111111;
20'b01100010000100100000: color_data = 12'b000011111111;
20'b01100010000100100100: color_data = 12'b000001101111;
20'b01100010000100100101: color_data = 12'b000001101111;
20'b01100010000100100110: color_data = 12'b000001101111;
20'b01100010000100100111: color_data = 12'b000001101111;
20'b01100010000100101000: color_data = 12'b000001101111;
20'b01100010000100101001: color_data = 12'b000001101111;
20'b01100010000100101010: color_data = 12'b000001101111;
20'b01100010000100101011: color_data = 12'b000001101111;
20'b01100010000100101100: color_data = 12'b000001101111;
20'b01100010000100101101: color_data = 12'b000001101111;
20'b01100010000100101110: color_data = 12'b000001101111;
20'b01100010000100101111: color_data = 12'b000001101111;
20'b01100010000100110000: color_data = 12'b000001101111;
20'b01100010000100110001: color_data = 12'b000001101111;
20'b01100010000100110010: color_data = 12'b000001101111;
20'b01100010000100110011: color_data = 12'b000001101111;
20'b01100010000100110100: color_data = 12'b000001101111;
20'b01100010000100110101: color_data = 12'b000001101111;
20'b01100010000100111001: color_data = 12'b000011110000;
20'b01100010000100111010: color_data = 12'b000011110000;
20'b01100010000100111011: color_data = 12'b000011110000;
20'b01100010000100111100: color_data = 12'b000011110000;
20'b01100010000100111101: color_data = 12'b000011110000;
20'b01100010000100111110: color_data = 12'b000011110000;
20'b01100010000100111111: color_data = 12'b000011110000;
20'b01100010000101000000: color_data = 12'b000011110000;
20'b01100010000101000001: color_data = 12'b000011110000;
20'b01100010000101000010: color_data = 12'b000011110000;
20'b01100010000101000011: color_data = 12'b000011110000;
20'b01100010000101000100: color_data = 12'b000011110000;
20'b01100010000101000101: color_data = 12'b000011110000;
20'b01100010000101000110: color_data = 12'b000011110000;
20'b01100010000101000111: color_data = 12'b000011110000;
20'b01100010000101001000: color_data = 12'b000011110000;
20'b01100010000101001001: color_data = 12'b000011110000;
20'b01100010000101001010: color_data = 12'b000011110000;
20'b01100010000101100011: color_data = 12'b111100001111;
20'b01100010000101100100: color_data = 12'b111100001111;
20'b01100010000101100101: color_data = 12'b111100001111;
20'b01100010000101100110: color_data = 12'b111100001111;
20'b01100010000101100111: color_data = 12'b111100001111;
20'b01100010000101101000: color_data = 12'b111100001111;
20'b01100010000101101001: color_data = 12'b111100001111;
20'b01100010000101101010: color_data = 12'b111100001111;
20'b01100010000101101011: color_data = 12'b111100001111;
20'b01100010000101101100: color_data = 12'b111100001111;
20'b01100010000101101101: color_data = 12'b111100001111;
20'b01100010000101101110: color_data = 12'b111100001111;
20'b01100010000101101111: color_data = 12'b111100001111;
20'b01100010000101110000: color_data = 12'b111100001111;
20'b01100010000101110001: color_data = 12'b111100001111;
20'b01100010000101110010: color_data = 12'b111100001111;
20'b01100010000101110011: color_data = 12'b111100001111;
20'b01100010000101110100: color_data = 12'b111100001111;
20'b01100010000110001101: color_data = 12'b111100000000;
20'b01100010000110001110: color_data = 12'b111100000000;
20'b01100010000110001111: color_data = 12'b111100000000;
20'b01100010000110010000: color_data = 12'b111100000000;
20'b01100010000110010001: color_data = 12'b111100000000;
20'b01100010000110010010: color_data = 12'b111100000000;
20'b01100010000110010011: color_data = 12'b111100000000;
20'b01100010000110010100: color_data = 12'b111100000000;
20'b01100010000110010101: color_data = 12'b111100000000;
20'b01100010000110010110: color_data = 12'b111100000000;
20'b01100010000110010111: color_data = 12'b111100000000;
20'b01100010000110011000: color_data = 12'b111100000000;
20'b01100010000110011001: color_data = 12'b111100000000;
20'b01100010000110011010: color_data = 12'b111100000000;
20'b01100010000110011011: color_data = 12'b111100000000;
20'b01100010000110011100: color_data = 12'b111100000000;
20'b01100010000110011101: color_data = 12'b111100000000;
20'b01100010000110011110: color_data = 12'b111100000000;
20'b01100010010011111010: color_data = 12'b000011111111;
20'b01100010010011111011: color_data = 12'b000011111111;
20'b01100010010011111100: color_data = 12'b000011111111;
20'b01100010010011111101: color_data = 12'b000011111111;
20'b01100010010011111110: color_data = 12'b000011111111;
20'b01100010010011111111: color_data = 12'b000011111111;
20'b01100010010100000000: color_data = 12'b000011111111;
20'b01100010010100000001: color_data = 12'b000011111111;
20'b01100010010100000010: color_data = 12'b000011111111;
20'b01100010010100000011: color_data = 12'b000011111111;
20'b01100010010100000100: color_data = 12'b000011111111;
20'b01100010010100000101: color_data = 12'b000011111111;
20'b01100010010100000110: color_data = 12'b000011111111;
20'b01100010010100000111: color_data = 12'b000011111111;
20'b01100010010100001000: color_data = 12'b000011111111;
20'b01100010010100001001: color_data = 12'b000011111111;
20'b01100010010100001010: color_data = 12'b000011111111;
20'b01100010010100001011: color_data = 12'b000011111111;
20'b01100010010100001111: color_data = 12'b000011111111;
20'b01100010010100010000: color_data = 12'b000011111111;
20'b01100010010100010001: color_data = 12'b000011111111;
20'b01100010010100010010: color_data = 12'b000011111111;
20'b01100010010100010011: color_data = 12'b000011111111;
20'b01100010010100010100: color_data = 12'b000011111111;
20'b01100010010100010101: color_data = 12'b000011111111;
20'b01100010010100010110: color_data = 12'b000011111111;
20'b01100010010100010111: color_data = 12'b000011111111;
20'b01100010010100011000: color_data = 12'b000011111111;
20'b01100010010100011001: color_data = 12'b000011111111;
20'b01100010010100011010: color_data = 12'b000011111111;
20'b01100010010100011011: color_data = 12'b000011111111;
20'b01100010010100011100: color_data = 12'b000011111111;
20'b01100010010100011101: color_data = 12'b000011111111;
20'b01100010010100011110: color_data = 12'b000011111111;
20'b01100010010100011111: color_data = 12'b000011111111;
20'b01100010010100100000: color_data = 12'b000011111111;
20'b01100010010100100100: color_data = 12'b000001101111;
20'b01100010010100100101: color_data = 12'b000001101111;
20'b01100010010100100110: color_data = 12'b000001101111;
20'b01100010010100100111: color_data = 12'b000001101111;
20'b01100010010100101000: color_data = 12'b000001101111;
20'b01100010010100101001: color_data = 12'b000001101111;
20'b01100010010100101010: color_data = 12'b000001101111;
20'b01100010010100101011: color_data = 12'b000001101111;
20'b01100010010100101100: color_data = 12'b000001101111;
20'b01100010010100101101: color_data = 12'b000001101111;
20'b01100010010100101110: color_data = 12'b000001101111;
20'b01100010010100101111: color_data = 12'b000001101111;
20'b01100010010100110000: color_data = 12'b000001101111;
20'b01100010010100110001: color_data = 12'b000001101111;
20'b01100010010100110010: color_data = 12'b000001101111;
20'b01100010010100110011: color_data = 12'b000001101111;
20'b01100010010100110100: color_data = 12'b000001101111;
20'b01100010010100110101: color_data = 12'b000001101111;
20'b01100010010100111001: color_data = 12'b000011110000;
20'b01100010010100111010: color_data = 12'b000011110000;
20'b01100010010100111011: color_data = 12'b000011110000;
20'b01100010010100111100: color_data = 12'b000011110000;
20'b01100010010100111101: color_data = 12'b000011110000;
20'b01100010010100111110: color_data = 12'b000011110000;
20'b01100010010100111111: color_data = 12'b000011110000;
20'b01100010010101000000: color_data = 12'b000011110000;
20'b01100010010101000001: color_data = 12'b000011110000;
20'b01100010010101000010: color_data = 12'b000011110000;
20'b01100010010101000011: color_data = 12'b000011110000;
20'b01100010010101000100: color_data = 12'b000011110000;
20'b01100010010101000101: color_data = 12'b000011110000;
20'b01100010010101000110: color_data = 12'b000011110000;
20'b01100010010101000111: color_data = 12'b000011110000;
20'b01100010010101001000: color_data = 12'b000011110000;
20'b01100010010101001001: color_data = 12'b000011110000;
20'b01100010010101001010: color_data = 12'b000011110000;
20'b01100010010101100011: color_data = 12'b111100001111;
20'b01100010010101100100: color_data = 12'b111100001111;
20'b01100010010101100101: color_data = 12'b111100001111;
20'b01100010010101100110: color_data = 12'b111100001111;
20'b01100010010101100111: color_data = 12'b111100001111;
20'b01100010010101101000: color_data = 12'b111100001111;
20'b01100010010101101001: color_data = 12'b111100001111;
20'b01100010010101101010: color_data = 12'b111100001111;
20'b01100010010101101011: color_data = 12'b111100001111;
20'b01100010010101101100: color_data = 12'b111100001111;
20'b01100010010101101101: color_data = 12'b111100001111;
20'b01100010010101101110: color_data = 12'b111100001111;
20'b01100010010101101111: color_data = 12'b111100001111;
20'b01100010010101110000: color_data = 12'b111100001111;
20'b01100010010101110001: color_data = 12'b111100001111;
20'b01100010010101110010: color_data = 12'b111100001111;
20'b01100010010101110011: color_data = 12'b111100001111;
20'b01100010010101110100: color_data = 12'b111100001111;
20'b01100010010110001101: color_data = 12'b111100000000;
20'b01100010010110001110: color_data = 12'b111100000000;
20'b01100010010110001111: color_data = 12'b111100000000;
20'b01100010010110010000: color_data = 12'b111100000000;
20'b01100010010110010001: color_data = 12'b111100000000;
20'b01100010010110010010: color_data = 12'b111100000000;
20'b01100010010110010011: color_data = 12'b111100000000;
20'b01100010010110010100: color_data = 12'b111100000000;
20'b01100010010110010101: color_data = 12'b111100000000;
20'b01100010010110010110: color_data = 12'b111100000000;
20'b01100010010110010111: color_data = 12'b111100000000;
20'b01100010010110011000: color_data = 12'b111100000000;
20'b01100010010110011001: color_data = 12'b111100000000;
20'b01100010010110011010: color_data = 12'b111100000000;
20'b01100010010110011011: color_data = 12'b111100000000;
20'b01100010010110011100: color_data = 12'b111100000000;
20'b01100010010110011101: color_data = 12'b111100000000;
20'b01100010010110011110: color_data = 12'b111100000000;
20'b01100010100011111010: color_data = 12'b000011111111;
20'b01100010100011111011: color_data = 12'b000011111111;
20'b01100010100011111100: color_data = 12'b000011111111;
20'b01100010100011111101: color_data = 12'b000011111111;
20'b01100010100011111110: color_data = 12'b000011111111;
20'b01100010100011111111: color_data = 12'b000011111111;
20'b01100010100100000000: color_data = 12'b000011111111;
20'b01100010100100000001: color_data = 12'b000011111111;
20'b01100010100100000010: color_data = 12'b000011111111;
20'b01100010100100000011: color_data = 12'b000011111111;
20'b01100010100100000100: color_data = 12'b000011111111;
20'b01100010100100000101: color_data = 12'b000011111111;
20'b01100010100100000110: color_data = 12'b000011111111;
20'b01100010100100000111: color_data = 12'b000011111111;
20'b01100010100100001000: color_data = 12'b000011111111;
20'b01100010100100001001: color_data = 12'b000011111111;
20'b01100010100100001010: color_data = 12'b000011111111;
20'b01100010100100001011: color_data = 12'b000011111111;
20'b01100010100100001111: color_data = 12'b000011111111;
20'b01100010100100010000: color_data = 12'b000011111111;
20'b01100010100100010001: color_data = 12'b000011111111;
20'b01100010100100010010: color_data = 12'b000011111111;
20'b01100010100100010011: color_data = 12'b000011111111;
20'b01100010100100010100: color_data = 12'b000011111111;
20'b01100010100100010101: color_data = 12'b000011111111;
20'b01100010100100010110: color_data = 12'b000011111111;
20'b01100010100100010111: color_data = 12'b000011111111;
20'b01100010100100011000: color_data = 12'b000011111111;
20'b01100010100100011001: color_data = 12'b000011111111;
20'b01100010100100011010: color_data = 12'b000011111111;
20'b01100010100100011011: color_data = 12'b000011111111;
20'b01100010100100011100: color_data = 12'b000011111111;
20'b01100010100100011101: color_data = 12'b000011111111;
20'b01100010100100011110: color_data = 12'b000011111111;
20'b01100010100100011111: color_data = 12'b000011111111;
20'b01100010100100100000: color_data = 12'b000011111111;
20'b01100010100100100100: color_data = 12'b000001101111;
20'b01100010100100100101: color_data = 12'b000001101111;
20'b01100010100100100110: color_data = 12'b000001101111;
20'b01100010100100100111: color_data = 12'b000001101111;
20'b01100010100100101000: color_data = 12'b000001101111;
20'b01100010100100101001: color_data = 12'b000001101111;
20'b01100010100100101010: color_data = 12'b000001101111;
20'b01100010100100101011: color_data = 12'b000001101111;
20'b01100010100100101100: color_data = 12'b000001101111;
20'b01100010100100101101: color_data = 12'b000001101111;
20'b01100010100100101110: color_data = 12'b000001101111;
20'b01100010100100101111: color_data = 12'b000001101111;
20'b01100010100100110000: color_data = 12'b000001101111;
20'b01100010100100110001: color_data = 12'b000001101111;
20'b01100010100100110010: color_data = 12'b000001101111;
20'b01100010100100110011: color_data = 12'b000001101111;
20'b01100010100100110100: color_data = 12'b000001101111;
20'b01100010100100110101: color_data = 12'b000001101111;
20'b01100010100100111001: color_data = 12'b000011110000;
20'b01100010100100111010: color_data = 12'b000011110000;
20'b01100010100100111011: color_data = 12'b000011110000;
20'b01100010100100111100: color_data = 12'b000011110000;
20'b01100010100100111101: color_data = 12'b000011110000;
20'b01100010100100111110: color_data = 12'b000011110000;
20'b01100010100100111111: color_data = 12'b000011110000;
20'b01100010100101000000: color_data = 12'b000011110000;
20'b01100010100101000001: color_data = 12'b000011110000;
20'b01100010100101000010: color_data = 12'b000011110000;
20'b01100010100101000011: color_data = 12'b000011110000;
20'b01100010100101000100: color_data = 12'b000011110000;
20'b01100010100101000101: color_data = 12'b000011110000;
20'b01100010100101000110: color_data = 12'b000011110000;
20'b01100010100101000111: color_data = 12'b000011110000;
20'b01100010100101001000: color_data = 12'b000011110000;
20'b01100010100101001001: color_data = 12'b000011110000;
20'b01100010100101001010: color_data = 12'b000011110000;
20'b01100010100101100011: color_data = 12'b111100001111;
20'b01100010100101100100: color_data = 12'b111100001111;
20'b01100010100101100101: color_data = 12'b111100001111;
20'b01100010100101100110: color_data = 12'b111100001111;
20'b01100010100101100111: color_data = 12'b111100001111;
20'b01100010100101101000: color_data = 12'b111100001111;
20'b01100010100101101001: color_data = 12'b111100001111;
20'b01100010100101101010: color_data = 12'b111100001111;
20'b01100010100101101011: color_data = 12'b111100001111;
20'b01100010100101101100: color_data = 12'b111100001111;
20'b01100010100101101101: color_data = 12'b111100001111;
20'b01100010100101101110: color_data = 12'b111100001111;
20'b01100010100101101111: color_data = 12'b111100001111;
20'b01100010100101110000: color_data = 12'b111100001111;
20'b01100010100101110001: color_data = 12'b111100001111;
20'b01100010100101110010: color_data = 12'b111100001111;
20'b01100010100101110011: color_data = 12'b111100001111;
20'b01100010100101110100: color_data = 12'b111100001111;
20'b01100010100110001101: color_data = 12'b111100000000;
20'b01100010100110001110: color_data = 12'b111100000000;
20'b01100010100110001111: color_data = 12'b111100000000;
20'b01100010100110010000: color_data = 12'b111100000000;
20'b01100010100110010001: color_data = 12'b111100000000;
20'b01100010100110010010: color_data = 12'b111100000000;
20'b01100010100110010011: color_data = 12'b111100000000;
20'b01100010100110010100: color_data = 12'b111100000000;
20'b01100010100110010101: color_data = 12'b111100000000;
20'b01100010100110010110: color_data = 12'b111100000000;
20'b01100010100110010111: color_data = 12'b111100000000;
20'b01100010100110011000: color_data = 12'b111100000000;
20'b01100010100110011001: color_data = 12'b111100000000;
20'b01100010100110011010: color_data = 12'b111100000000;
20'b01100010100110011011: color_data = 12'b111100000000;
20'b01100010100110011100: color_data = 12'b111100000000;
20'b01100010100110011101: color_data = 12'b111100000000;
20'b01100010100110011110: color_data = 12'b111100000000;
20'b01100010110011111010: color_data = 12'b000011111111;
20'b01100010110011111011: color_data = 12'b000011111111;
20'b01100010110011111100: color_data = 12'b000011111111;
20'b01100010110011111101: color_data = 12'b000011111111;
20'b01100010110011111110: color_data = 12'b000011111111;
20'b01100010110011111111: color_data = 12'b000011111111;
20'b01100010110100000000: color_data = 12'b000011111111;
20'b01100010110100000001: color_data = 12'b000011111111;
20'b01100010110100000010: color_data = 12'b000011111111;
20'b01100010110100000011: color_data = 12'b000011111111;
20'b01100010110100000100: color_data = 12'b000011111111;
20'b01100010110100000101: color_data = 12'b000011111111;
20'b01100010110100000110: color_data = 12'b000011111111;
20'b01100010110100000111: color_data = 12'b000011111111;
20'b01100010110100001000: color_data = 12'b000011111111;
20'b01100010110100001001: color_data = 12'b000011111111;
20'b01100010110100001010: color_data = 12'b000011111111;
20'b01100010110100001011: color_data = 12'b000011111111;
20'b01100010110100001111: color_data = 12'b000011111111;
20'b01100010110100010000: color_data = 12'b000011111111;
20'b01100010110100010001: color_data = 12'b000011111111;
20'b01100010110100010010: color_data = 12'b000011111111;
20'b01100010110100010011: color_data = 12'b000011111111;
20'b01100010110100010100: color_data = 12'b000011111111;
20'b01100010110100010101: color_data = 12'b000011111111;
20'b01100010110100010110: color_data = 12'b000011111111;
20'b01100010110100010111: color_data = 12'b000011111111;
20'b01100010110100011000: color_data = 12'b000011111111;
20'b01100010110100011001: color_data = 12'b000011111111;
20'b01100010110100011010: color_data = 12'b000011111111;
20'b01100010110100011011: color_data = 12'b000011111111;
20'b01100010110100011100: color_data = 12'b000011111111;
20'b01100010110100011101: color_data = 12'b000011111111;
20'b01100010110100011110: color_data = 12'b000011111111;
20'b01100010110100011111: color_data = 12'b000011111111;
20'b01100010110100100000: color_data = 12'b000011111111;
20'b01100010110100100100: color_data = 12'b000001101111;
20'b01100010110100100101: color_data = 12'b000001101111;
20'b01100010110100100110: color_data = 12'b000001101111;
20'b01100010110100100111: color_data = 12'b000001101111;
20'b01100010110100101000: color_data = 12'b000001101111;
20'b01100010110100101001: color_data = 12'b000001101111;
20'b01100010110100101010: color_data = 12'b000001101111;
20'b01100010110100101011: color_data = 12'b000001101111;
20'b01100010110100101100: color_data = 12'b000001101111;
20'b01100010110100101101: color_data = 12'b000001101111;
20'b01100010110100101110: color_data = 12'b000001101111;
20'b01100010110100101111: color_data = 12'b000001101111;
20'b01100010110100110000: color_data = 12'b000001101111;
20'b01100010110100110001: color_data = 12'b000001101111;
20'b01100010110100110010: color_data = 12'b000001101111;
20'b01100010110100110011: color_data = 12'b000001101111;
20'b01100010110100110100: color_data = 12'b000001101111;
20'b01100010110100110101: color_data = 12'b000001101111;
20'b01100010110100111001: color_data = 12'b000011110000;
20'b01100010110100111010: color_data = 12'b000011110000;
20'b01100010110100111011: color_data = 12'b000011110000;
20'b01100010110100111100: color_data = 12'b000011110000;
20'b01100010110100111101: color_data = 12'b000011110000;
20'b01100010110100111110: color_data = 12'b000011110000;
20'b01100010110100111111: color_data = 12'b000011110000;
20'b01100010110101000000: color_data = 12'b000011110000;
20'b01100010110101000001: color_data = 12'b000011110000;
20'b01100010110101000010: color_data = 12'b000011110000;
20'b01100010110101000011: color_data = 12'b000011110000;
20'b01100010110101000100: color_data = 12'b000011110000;
20'b01100010110101000101: color_data = 12'b000011110000;
20'b01100010110101000110: color_data = 12'b000011110000;
20'b01100010110101000111: color_data = 12'b000011110000;
20'b01100010110101001000: color_data = 12'b000011110000;
20'b01100010110101001001: color_data = 12'b000011110000;
20'b01100010110101001010: color_data = 12'b000011110000;
20'b01100010110101100011: color_data = 12'b111100001111;
20'b01100010110101100100: color_data = 12'b111100001111;
20'b01100010110101100101: color_data = 12'b111100001111;
20'b01100010110101100110: color_data = 12'b111100001111;
20'b01100010110101100111: color_data = 12'b111100001111;
20'b01100010110101101000: color_data = 12'b111100001111;
20'b01100010110101101001: color_data = 12'b111100001111;
20'b01100010110101101010: color_data = 12'b111100001111;
20'b01100010110101101011: color_data = 12'b111100001111;
20'b01100010110101101100: color_data = 12'b111100001111;
20'b01100010110101101101: color_data = 12'b111100001111;
20'b01100010110101101110: color_data = 12'b111100001111;
20'b01100010110101101111: color_data = 12'b111100001111;
20'b01100010110101110000: color_data = 12'b111100001111;
20'b01100010110101110001: color_data = 12'b111100001111;
20'b01100010110101110010: color_data = 12'b111100001111;
20'b01100010110101110011: color_data = 12'b111100001111;
20'b01100010110101110100: color_data = 12'b111100001111;
20'b01100010110110001101: color_data = 12'b111100000000;
20'b01100010110110001110: color_data = 12'b111100000000;
20'b01100010110110001111: color_data = 12'b111100000000;
20'b01100010110110010000: color_data = 12'b111100000000;
20'b01100010110110010001: color_data = 12'b111100000000;
20'b01100010110110010010: color_data = 12'b111100000000;
20'b01100010110110010011: color_data = 12'b111100000000;
20'b01100010110110010100: color_data = 12'b111100000000;
20'b01100010110110010101: color_data = 12'b111100000000;
20'b01100010110110010110: color_data = 12'b111100000000;
20'b01100010110110010111: color_data = 12'b111100000000;
20'b01100010110110011000: color_data = 12'b111100000000;
20'b01100010110110011001: color_data = 12'b111100000000;
20'b01100010110110011010: color_data = 12'b111100000000;
20'b01100010110110011011: color_data = 12'b111100000000;
20'b01100010110110011100: color_data = 12'b111100000000;
20'b01100010110110011101: color_data = 12'b111100000000;
20'b01100010110110011110: color_data = 12'b111100000000;
20'b01100011000011111010: color_data = 12'b000011111111;
20'b01100011000011111011: color_data = 12'b000011111111;
20'b01100011000011111100: color_data = 12'b000011111111;
20'b01100011000011111101: color_data = 12'b000011111111;
20'b01100011000011111110: color_data = 12'b000011111111;
20'b01100011000011111111: color_data = 12'b000011111111;
20'b01100011000100000000: color_data = 12'b000011111111;
20'b01100011000100000001: color_data = 12'b000011111111;
20'b01100011000100000010: color_data = 12'b000011111111;
20'b01100011000100000011: color_data = 12'b000011111111;
20'b01100011000100000100: color_data = 12'b000011111111;
20'b01100011000100000101: color_data = 12'b000011111111;
20'b01100011000100000110: color_data = 12'b000011111111;
20'b01100011000100000111: color_data = 12'b000011111111;
20'b01100011000100001000: color_data = 12'b000011111111;
20'b01100011000100001001: color_data = 12'b000011111111;
20'b01100011000100001010: color_data = 12'b000011111111;
20'b01100011000100001011: color_data = 12'b000011111111;
20'b01100011000100001111: color_data = 12'b000011111111;
20'b01100011000100010000: color_data = 12'b000011111111;
20'b01100011000100010001: color_data = 12'b000011111111;
20'b01100011000100010010: color_data = 12'b000011111111;
20'b01100011000100010011: color_data = 12'b000011111111;
20'b01100011000100010100: color_data = 12'b000011111111;
20'b01100011000100010101: color_data = 12'b000011111111;
20'b01100011000100010110: color_data = 12'b000011111111;
20'b01100011000100010111: color_data = 12'b000011111111;
20'b01100011000100011000: color_data = 12'b000011111111;
20'b01100011000100011001: color_data = 12'b000011111111;
20'b01100011000100011010: color_data = 12'b000011111111;
20'b01100011000100011011: color_data = 12'b000011111111;
20'b01100011000100011100: color_data = 12'b000011111111;
20'b01100011000100011101: color_data = 12'b000011111111;
20'b01100011000100011110: color_data = 12'b000011111111;
20'b01100011000100011111: color_data = 12'b000011111111;
20'b01100011000100100000: color_data = 12'b000011111111;
20'b01100011000100100100: color_data = 12'b000001101111;
20'b01100011000100100101: color_data = 12'b000001101111;
20'b01100011000100100110: color_data = 12'b000001101111;
20'b01100011000100100111: color_data = 12'b000001101111;
20'b01100011000100101000: color_data = 12'b000001101111;
20'b01100011000100101001: color_data = 12'b000001101111;
20'b01100011000100101010: color_data = 12'b000001101111;
20'b01100011000100101011: color_data = 12'b000001101111;
20'b01100011000100101100: color_data = 12'b000001101111;
20'b01100011000100101101: color_data = 12'b000001101111;
20'b01100011000100101110: color_data = 12'b000001101111;
20'b01100011000100101111: color_data = 12'b000001101111;
20'b01100011000100110000: color_data = 12'b000001101111;
20'b01100011000100110001: color_data = 12'b000001101111;
20'b01100011000100110010: color_data = 12'b000001101111;
20'b01100011000100110011: color_data = 12'b000001101111;
20'b01100011000100110100: color_data = 12'b000001101111;
20'b01100011000100110101: color_data = 12'b000001101111;
20'b01100011000100111001: color_data = 12'b000011110000;
20'b01100011000100111010: color_data = 12'b000011110000;
20'b01100011000100111011: color_data = 12'b000011110000;
20'b01100011000100111100: color_data = 12'b000011110000;
20'b01100011000100111101: color_data = 12'b000011110000;
20'b01100011000100111110: color_data = 12'b000011110000;
20'b01100011000100111111: color_data = 12'b000011110000;
20'b01100011000101000000: color_data = 12'b000011110000;
20'b01100011000101000001: color_data = 12'b000011110000;
20'b01100011000101000010: color_data = 12'b000011110000;
20'b01100011000101000011: color_data = 12'b000011110000;
20'b01100011000101000100: color_data = 12'b000011110000;
20'b01100011000101000101: color_data = 12'b000011110000;
20'b01100011000101000110: color_data = 12'b000011110000;
20'b01100011000101000111: color_data = 12'b000011110000;
20'b01100011000101001000: color_data = 12'b000011110000;
20'b01100011000101001001: color_data = 12'b000011110000;
20'b01100011000101001010: color_data = 12'b000011110000;
20'b01100011000101100011: color_data = 12'b111100001111;
20'b01100011000101100100: color_data = 12'b111100001111;
20'b01100011000101100101: color_data = 12'b111100001111;
20'b01100011000101100110: color_data = 12'b111100001111;
20'b01100011000101100111: color_data = 12'b111100001111;
20'b01100011000101101000: color_data = 12'b111100001111;
20'b01100011000101101001: color_data = 12'b111100001111;
20'b01100011000101101010: color_data = 12'b111100001111;
20'b01100011000101101011: color_data = 12'b111100001111;
20'b01100011000101101100: color_data = 12'b111100001111;
20'b01100011000101101101: color_data = 12'b111100001111;
20'b01100011000101101110: color_data = 12'b111100001111;
20'b01100011000101101111: color_data = 12'b111100001111;
20'b01100011000101110000: color_data = 12'b111100001111;
20'b01100011000101110001: color_data = 12'b111100001111;
20'b01100011000101110010: color_data = 12'b111100001111;
20'b01100011000101110011: color_data = 12'b111100001111;
20'b01100011000101110100: color_data = 12'b111100001111;
20'b01100011000110001101: color_data = 12'b111100000000;
20'b01100011000110001110: color_data = 12'b111100000000;
20'b01100011000110001111: color_data = 12'b111100000000;
20'b01100011000110010000: color_data = 12'b111100000000;
20'b01100011000110010001: color_data = 12'b111100000000;
20'b01100011000110010010: color_data = 12'b111100000000;
20'b01100011000110010011: color_data = 12'b111100000000;
20'b01100011000110010100: color_data = 12'b111100000000;
20'b01100011000110010101: color_data = 12'b111100000000;
20'b01100011000110010110: color_data = 12'b111100000000;
20'b01100011000110010111: color_data = 12'b111100000000;
20'b01100011000110011000: color_data = 12'b111100000000;
20'b01100011000110011001: color_data = 12'b111100000000;
20'b01100011000110011010: color_data = 12'b111100000000;
20'b01100011000110011011: color_data = 12'b111100000000;
20'b01100011000110011100: color_data = 12'b111100000000;
20'b01100011000110011101: color_data = 12'b111100000000;
20'b01100011000110011110: color_data = 12'b111100000000;
20'b01100100000011111010: color_data = 12'b000001101111;
20'b01100100000011111011: color_data = 12'b000001101111;
20'b01100100000011111100: color_data = 12'b000001101111;
20'b01100100000011111101: color_data = 12'b000001101111;
20'b01100100000011111110: color_data = 12'b000001101111;
20'b01100100000011111111: color_data = 12'b000001101111;
20'b01100100000100000000: color_data = 12'b000001101111;
20'b01100100000100000001: color_data = 12'b000001101111;
20'b01100100000100000010: color_data = 12'b000001101111;
20'b01100100000100000011: color_data = 12'b000001101111;
20'b01100100000100000100: color_data = 12'b000001101111;
20'b01100100000100000101: color_data = 12'b000001101111;
20'b01100100000100000110: color_data = 12'b000001101111;
20'b01100100000100000111: color_data = 12'b000001101111;
20'b01100100000100001000: color_data = 12'b000001101111;
20'b01100100000100001001: color_data = 12'b000001101111;
20'b01100100000100001010: color_data = 12'b000001101111;
20'b01100100000100001011: color_data = 12'b000001101111;
20'b01100100000100001111: color_data = 12'b000001101111;
20'b01100100000100010000: color_data = 12'b000001101111;
20'b01100100000100010001: color_data = 12'b000001101111;
20'b01100100000100010010: color_data = 12'b000001101111;
20'b01100100000100010011: color_data = 12'b000001101111;
20'b01100100000100010100: color_data = 12'b000001101111;
20'b01100100000100010101: color_data = 12'b000001101111;
20'b01100100000100010110: color_data = 12'b000001101111;
20'b01100100000100010111: color_data = 12'b000001101111;
20'b01100100000100011000: color_data = 12'b000001101111;
20'b01100100000100011001: color_data = 12'b000001101111;
20'b01100100000100011010: color_data = 12'b000001101111;
20'b01100100000100011011: color_data = 12'b000001101111;
20'b01100100000100011100: color_data = 12'b000001101111;
20'b01100100000100011101: color_data = 12'b000001101111;
20'b01100100000100011110: color_data = 12'b000001101111;
20'b01100100000100011111: color_data = 12'b000001101111;
20'b01100100000100100000: color_data = 12'b000001101111;
20'b01100100000100100100: color_data = 12'b000001101111;
20'b01100100000100100101: color_data = 12'b000001101111;
20'b01100100000100100110: color_data = 12'b000001101111;
20'b01100100000100100111: color_data = 12'b000001101111;
20'b01100100000100101000: color_data = 12'b000001101111;
20'b01100100000100101001: color_data = 12'b000001101111;
20'b01100100000100101010: color_data = 12'b000001101111;
20'b01100100000100101011: color_data = 12'b000001101111;
20'b01100100000100101100: color_data = 12'b000001101111;
20'b01100100000100101101: color_data = 12'b000001101111;
20'b01100100000100101110: color_data = 12'b000001101111;
20'b01100100000100101111: color_data = 12'b000001101111;
20'b01100100000100110000: color_data = 12'b000001101111;
20'b01100100000100110001: color_data = 12'b000001101111;
20'b01100100000100110010: color_data = 12'b000001101111;
20'b01100100000100110011: color_data = 12'b000001101111;
20'b01100100000100110100: color_data = 12'b000001101111;
20'b01100100000100110101: color_data = 12'b000001101111;
20'b01100100000100111001: color_data = 12'b000011110000;
20'b01100100000100111010: color_data = 12'b000011110000;
20'b01100100000100111011: color_data = 12'b000011110000;
20'b01100100000100111100: color_data = 12'b000011110000;
20'b01100100000100111101: color_data = 12'b000011110000;
20'b01100100000100111110: color_data = 12'b000011110000;
20'b01100100000100111111: color_data = 12'b000011110000;
20'b01100100000101000000: color_data = 12'b000011110000;
20'b01100100000101000001: color_data = 12'b000011110000;
20'b01100100000101000010: color_data = 12'b000011110000;
20'b01100100000101000011: color_data = 12'b000011110000;
20'b01100100000101000100: color_data = 12'b000011110000;
20'b01100100000101000101: color_data = 12'b000011110000;
20'b01100100000101000110: color_data = 12'b000011110000;
20'b01100100000101000111: color_data = 12'b000011110000;
20'b01100100000101001000: color_data = 12'b000011110000;
20'b01100100000101001001: color_data = 12'b000011110000;
20'b01100100000101001010: color_data = 12'b000011110000;
20'b01100100000101001110: color_data = 12'b000011110000;
20'b01100100000101001111: color_data = 12'b000011110000;
20'b01100100000101010000: color_data = 12'b000011110000;
20'b01100100000101010001: color_data = 12'b000011110000;
20'b01100100000101010010: color_data = 12'b000011110000;
20'b01100100000101010011: color_data = 12'b000011110000;
20'b01100100000101010100: color_data = 12'b000011110000;
20'b01100100000101010101: color_data = 12'b000011110000;
20'b01100100000101010110: color_data = 12'b000011110000;
20'b01100100000101010111: color_data = 12'b000011110000;
20'b01100100000101011000: color_data = 12'b000011110000;
20'b01100100000101011001: color_data = 12'b000011110000;
20'b01100100000101011010: color_data = 12'b000011110000;
20'b01100100000101011011: color_data = 12'b000011110000;
20'b01100100000101011100: color_data = 12'b000011110000;
20'b01100100000101011101: color_data = 12'b000011110000;
20'b01100100000101011110: color_data = 12'b000011110000;
20'b01100100000101011111: color_data = 12'b000011110000;
20'b01100100000101100011: color_data = 12'b111100001111;
20'b01100100000101100100: color_data = 12'b111100001111;
20'b01100100000101100101: color_data = 12'b111100001111;
20'b01100100000101100110: color_data = 12'b111100001111;
20'b01100100000101100111: color_data = 12'b111100001111;
20'b01100100000101101000: color_data = 12'b111100001111;
20'b01100100000101101001: color_data = 12'b111100001111;
20'b01100100000101101010: color_data = 12'b111100001111;
20'b01100100000101101011: color_data = 12'b111100001111;
20'b01100100000101101100: color_data = 12'b111100001111;
20'b01100100000101101101: color_data = 12'b111100001111;
20'b01100100000101101110: color_data = 12'b111100001111;
20'b01100100000101101111: color_data = 12'b111100001111;
20'b01100100000101110000: color_data = 12'b111100001111;
20'b01100100000101110001: color_data = 12'b111100001111;
20'b01100100000101110010: color_data = 12'b111100001111;
20'b01100100000101110011: color_data = 12'b111100001111;
20'b01100100000101110100: color_data = 12'b111100001111;
20'b01100100000101111000: color_data = 12'b111100001111;
20'b01100100000101111001: color_data = 12'b111100001111;
20'b01100100000101111010: color_data = 12'b111100001111;
20'b01100100000101111011: color_data = 12'b111100001111;
20'b01100100000101111100: color_data = 12'b111100001111;
20'b01100100000101111101: color_data = 12'b111100001111;
20'b01100100000101111110: color_data = 12'b111100001111;
20'b01100100000101111111: color_data = 12'b111100001111;
20'b01100100000110000000: color_data = 12'b111100001111;
20'b01100100000110000001: color_data = 12'b111100001111;
20'b01100100000110000010: color_data = 12'b111100001111;
20'b01100100000110000011: color_data = 12'b111100001111;
20'b01100100000110000100: color_data = 12'b111100001111;
20'b01100100000110000101: color_data = 12'b111100001111;
20'b01100100000110000110: color_data = 12'b111100001111;
20'b01100100000110000111: color_data = 12'b111100001111;
20'b01100100000110001000: color_data = 12'b111100001111;
20'b01100100000110001001: color_data = 12'b111100001111;
20'b01100100000110001101: color_data = 12'b111100000000;
20'b01100100000110001110: color_data = 12'b111100000000;
20'b01100100000110001111: color_data = 12'b111100000000;
20'b01100100000110010000: color_data = 12'b111100000000;
20'b01100100000110010001: color_data = 12'b111100000000;
20'b01100100000110010010: color_data = 12'b111100000000;
20'b01100100000110010011: color_data = 12'b111100000000;
20'b01100100000110010100: color_data = 12'b111100000000;
20'b01100100000110010101: color_data = 12'b111100000000;
20'b01100100000110010110: color_data = 12'b111100000000;
20'b01100100000110010111: color_data = 12'b111100000000;
20'b01100100000110011000: color_data = 12'b111100000000;
20'b01100100000110011001: color_data = 12'b111100000000;
20'b01100100000110011010: color_data = 12'b111100000000;
20'b01100100000110011011: color_data = 12'b111100000000;
20'b01100100000110011100: color_data = 12'b111100000000;
20'b01100100000110011101: color_data = 12'b111100000000;
20'b01100100000110011110: color_data = 12'b111100000000;
20'b01100100010011111010: color_data = 12'b000001101111;
20'b01100100010011111011: color_data = 12'b000001101111;
20'b01100100010011111100: color_data = 12'b000001101111;
20'b01100100010011111101: color_data = 12'b000001101111;
20'b01100100010011111110: color_data = 12'b000001101111;
20'b01100100010011111111: color_data = 12'b000001101111;
20'b01100100010100000000: color_data = 12'b000001101111;
20'b01100100010100000001: color_data = 12'b000001101111;
20'b01100100010100000010: color_data = 12'b000001101111;
20'b01100100010100000011: color_data = 12'b000001101111;
20'b01100100010100000100: color_data = 12'b000001101111;
20'b01100100010100000101: color_data = 12'b000001101111;
20'b01100100010100000110: color_data = 12'b000001101111;
20'b01100100010100000111: color_data = 12'b000001101111;
20'b01100100010100001000: color_data = 12'b000001101111;
20'b01100100010100001001: color_data = 12'b000001101111;
20'b01100100010100001010: color_data = 12'b000001101111;
20'b01100100010100001011: color_data = 12'b000001101111;
20'b01100100010100001111: color_data = 12'b000001101111;
20'b01100100010100010000: color_data = 12'b000001101111;
20'b01100100010100010001: color_data = 12'b000001101111;
20'b01100100010100010010: color_data = 12'b000001101111;
20'b01100100010100010011: color_data = 12'b000001101111;
20'b01100100010100010100: color_data = 12'b000001101111;
20'b01100100010100010101: color_data = 12'b000001101111;
20'b01100100010100010110: color_data = 12'b000001101111;
20'b01100100010100010111: color_data = 12'b000001101111;
20'b01100100010100011000: color_data = 12'b000001101111;
20'b01100100010100011001: color_data = 12'b000001101111;
20'b01100100010100011010: color_data = 12'b000001101111;
20'b01100100010100011011: color_data = 12'b000001101111;
20'b01100100010100011100: color_data = 12'b000001101111;
20'b01100100010100011101: color_data = 12'b000001101111;
20'b01100100010100011110: color_data = 12'b000001101111;
20'b01100100010100011111: color_data = 12'b000001101111;
20'b01100100010100100000: color_data = 12'b000001101111;
20'b01100100010100100100: color_data = 12'b000001101111;
20'b01100100010100100101: color_data = 12'b000001101111;
20'b01100100010100100110: color_data = 12'b000001101111;
20'b01100100010100100111: color_data = 12'b000001101111;
20'b01100100010100101000: color_data = 12'b000001101111;
20'b01100100010100101001: color_data = 12'b000001101111;
20'b01100100010100101010: color_data = 12'b000001101111;
20'b01100100010100101011: color_data = 12'b000001101111;
20'b01100100010100101100: color_data = 12'b000001101111;
20'b01100100010100101101: color_data = 12'b000001101111;
20'b01100100010100101110: color_data = 12'b000001101111;
20'b01100100010100101111: color_data = 12'b000001101111;
20'b01100100010100110000: color_data = 12'b000001101111;
20'b01100100010100110001: color_data = 12'b000001101111;
20'b01100100010100110010: color_data = 12'b000001101111;
20'b01100100010100110011: color_data = 12'b000001101111;
20'b01100100010100110100: color_data = 12'b000001101111;
20'b01100100010100110101: color_data = 12'b000001101111;
20'b01100100010100111001: color_data = 12'b000011110000;
20'b01100100010100111010: color_data = 12'b000011110000;
20'b01100100010100111011: color_data = 12'b000011110000;
20'b01100100010100111100: color_data = 12'b000011110000;
20'b01100100010100111101: color_data = 12'b000011110000;
20'b01100100010100111110: color_data = 12'b000011110000;
20'b01100100010100111111: color_data = 12'b000011110000;
20'b01100100010101000000: color_data = 12'b000011110000;
20'b01100100010101000001: color_data = 12'b000011110000;
20'b01100100010101000010: color_data = 12'b000011110000;
20'b01100100010101000011: color_data = 12'b000011110000;
20'b01100100010101000100: color_data = 12'b000011110000;
20'b01100100010101000101: color_data = 12'b000011110000;
20'b01100100010101000110: color_data = 12'b000011110000;
20'b01100100010101000111: color_data = 12'b000011110000;
20'b01100100010101001000: color_data = 12'b000011110000;
20'b01100100010101001001: color_data = 12'b000011110000;
20'b01100100010101001010: color_data = 12'b000011110000;
20'b01100100010101001110: color_data = 12'b000011110000;
20'b01100100010101001111: color_data = 12'b000011110000;
20'b01100100010101010000: color_data = 12'b000011110000;
20'b01100100010101010001: color_data = 12'b000011110000;
20'b01100100010101010010: color_data = 12'b000011110000;
20'b01100100010101010011: color_data = 12'b000011110000;
20'b01100100010101010100: color_data = 12'b000011110000;
20'b01100100010101010101: color_data = 12'b000011110000;
20'b01100100010101010110: color_data = 12'b000011110000;
20'b01100100010101010111: color_data = 12'b000011110000;
20'b01100100010101011000: color_data = 12'b000011110000;
20'b01100100010101011001: color_data = 12'b000011110000;
20'b01100100010101011010: color_data = 12'b000011110000;
20'b01100100010101011011: color_data = 12'b000011110000;
20'b01100100010101011100: color_data = 12'b000011110000;
20'b01100100010101011101: color_data = 12'b000011110000;
20'b01100100010101011110: color_data = 12'b000011110000;
20'b01100100010101011111: color_data = 12'b000011110000;
20'b01100100010101100011: color_data = 12'b111100001111;
20'b01100100010101100100: color_data = 12'b111100001111;
20'b01100100010101100101: color_data = 12'b111100001111;
20'b01100100010101100110: color_data = 12'b111100001111;
20'b01100100010101100111: color_data = 12'b111100001111;
20'b01100100010101101000: color_data = 12'b111100001111;
20'b01100100010101101001: color_data = 12'b111100001111;
20'b01100100010101101010: color_data = 12'b111100001111;
20'b01100100010101101011: color_data = 12'b111100001111;
20'b01100100010101101100: color_data = 12'b111100001111;
20'b01100100010101101101: color_data = 12'b111100001111;
20'b01100100010101101110: color_data = 12'b111100001111;
20'b01100100010101101111: color_data = 12'b111100001111;
20'b01100100010101110000: color_data = 12'b111100001111;
20'b01100100010101110001: color_data = 12'b111100001111;
20'b01100100010101110010: color_data = 12'b111100001111;
20'b01100100010101110011: color_data = 12'b111100001111;
20'b01100100010101110100: color_data = 12'b111100001111;
20'b01100100010101111000: color_data = 12'b111100001111;
20'b01100100010101111001: color_data = 12'b111100001111;
20'b01100100010101111010: color_data = 12'b111100001111;
20'b01100100010101111011: color_data = 12'b111100001111;
20'b01100100010101111100: color_data = 12'b111100001111;
20'b01100100010101111101: color_data = 12'b111100001111;
20'b01100100010101111110: color_data = 12'b111100001111;
20'b01100100010101111111: color_data = 12'b111100001111;
20'b01100100010110000000: color_data = 12'b111100001111;
20'b01100100010110000001: color_data = 12'b111100001111;
20'b01100100010110000010: color_data = 12'b111100001111;
20'b01100100010110000011: color_data = 12'b111100001111;
20'b01100100010110000100: color_data = 12'b111100001111;
20'b01100100010110000101: color_data = 12'b111100001111;
20'b01100100010110000110: color_data = 12'b111100001111;
20'b01100100010110000111: color_data = 12'b111100001111;
20'b01100100010110001000: color_data = 12'b111100001111;
20'b01100100010110001001: color_data = 12'b111100001111;
20'b01100100010110001101: color_data = 12'b111100000000;
20'b01100100010110001110: color_data = 12'b111100000000;
20'b01100100010110001111: color_data = 12'b111100000000;
20'b01100100010110010000: color_data = 12'b111100000000;
20'b01100100010110010001: color_data = 12'b111100000000;
20'b01100100010110010010: color_data = 12'b111100000000;
20'b01100100010110010011: color_data = 12'b111100000000;
20'b01100100010110010100: color_data = 12'b111100000000;
20'b01100100010110010101: color_data = 12'b111100000000;
20'b01100100010110010110: color_data = 12'b111100000000;
20'b01100100010110010111: color_data = 12'b111100000000;
20'b01100100010110011000: color_data = 12'b111100000000;
20'b01100100010110011001: color_data = 12'b111100000000;
20'b01100100010110011010: color_data = 12'b111100000000;
20'b01100100010110011011: color_data = 12'b111100000000;
20'b01100100010110011100: color_data = 12'b111100000000;
20'b01100100010110011101: color_data = 12'b111100000000;
20'b01100100010110011110: color_data = 12'b111100000000;
20'b01100100100011111010: color_data = 12'b000001101111;
20'b01100100100011111011: color_data = 12'b000001101111;
20'b01100100100011111100: color_data = 12'b000001101111;
20'b01100100100011111101: color_data = 12'b000001101111;
20'b01100100100011111110: color_data = 12'b000001101111;
20'b01100100100011111111: color_data = 12'b000001101111;
20'b01100100100100000000: color_data = 12'b000001101111;
20'b01100100100100000001: color_data = 12'b000001101111;
20'b01100100100100000010: color_data = 12'b000001101111;
20'b01100100100100000011: color_data = 12'b000001101111;
20'b01100100100100000100: color_data = 12'b000001101111;
20'b01100100100100000101: color_data = 12'b000001101111;
20'b01100100100100000110: color_data = 12'b000001101111;
20'b01100100100100000111: color_data = 12'b000001101111;
20'b01100100100100001000: color_data = 12'b000001101111;
20'b01100100100100001001: color_data = 12'b000001101111;
20'b01100100100100001010: color_data = 12'b000001101111;
20'b01100100100100001011: color_data = 12'b000001101111;
20'b01100100100100001111: color_data = 12'b000001101111;
20'b01100100100100010000: color_data = 12'b000001101111;
20'b01100100100100010001: color_data = 12'b000001101111;
20'b01100100100100010010: color_data = 12'b000001101111;
20'b01100100100100010011: color_data = 12'b000001101111;
20'b01100100100100010100: color_data = 12'b000001101111;
20'b01100100100100010101: color_data = 12'b000001101111;
20'b01100100100100010110: color_data = 12'b000001101111;
20'b01100100100100010111: color_data = 12'b000001101111;
20'b01100100100100011000: color_data = 12'b000001101111;
20'b01100100100100011001: color_data = 12'b000001101111;
20'b01100100100100011010: color_data = 12'b000001101111;
20'b01100100100100011011: color_data = 12'b000001101111;
20'b01100100100100011100: color_data = 12'b000001101111;
20'b01100100100100011101: color_data = 12'b000001101111;
20'b01100100100100011110: color_data = 12'b000001101111;
20'b01100100100100011111: color_data = 12'b000001101111;
20'b01100100100100100000: color_data = 12'b000001101111;
20'b01100100100100100100: color_data = 12'b000001101111;
20'b01100100100100100101: color_data = 12'b000001101111;
20'b01100100100100100110: color_data = 12'b000001101111;
20'b01100100100100100111: color_data = 12'b000001101111;
20'b01100100100100101000: color_data = 12'b000001101111;
20'b01100100100100101001: color_data = 12'b000001101111;
20'b01100100100100101010: color_data = 12'b000001101111;
20'b01100100100100101011: color_data = 12'b000001101111;
20'b01100100100100101100: color_data = 12'b000001101111;
20'b01100100100100101101: color_data = 12'b000001101111;
20'b01100100100100101110: color_data = 12'b000001101111;
20'b01100100100100101111: color_data = 12'b000001101111;
20'b01100100100100110000: color_data = 12'b000001101111;
20'b01100100100100110001: color_data = 12'b000001101111;
20'b01100100100100110010: color_data = 12'b000001101111;
20'b01100100100100110011: color_data = 12'b000001101111;
20'b01100100100100110100: color_data = 12'b000001101111;
20'b01100100100100110101: color_data = 12'b000001101111;
20'b01100100100100111001: color_data = 12'b000011110000;
20'b01100100100100111010: color_data = 12'b000011110000;
20'b01100100100100111011: color_data = 12'b000011110000;
20'b01100100100100111100: color_data = 12'b000011110000;
20'b01100100100100111101: color_data = 12'b000011110000;
20'b01100100100100111110: color_data = 12'b000011110000;
20'b01100100100100111111: color_data = 12'b000011110000;
20'b01100100100101000000: color_data = 12'b000011110000;
20'b01100100100101000001: color_data = 12'b000011110000;
20'b01100100100101000010: color_data = 12'b000011110000;
20'b01100100100101000011: color_data = 12'b000011110000;
20'b01100100100101000100: color_data = 12'b000011110000;
20'b01100100100101000101: color_data = 12'b000011110000;
20'b01100100100101000110: color_data = 12'b000011110000;
20'b01100100100101000111: color_data = 12'b000011110000;
20'b01100100100101001000: color_data = 12'b000011110000;
20'b01100100100101001001: color_data = 12'b000011110000;
20'b01100100100101001010: color_data = 12'b000011110000;
20'b01100100100101001110: color_data = 12'b000011110000;
20'b01100100100101001111: color_data = 12'b000011110000;
20'b01100100100101010000: color_data = 12'b000011110000;
20'b01100100100101010001: color_data = 12'b000011110000;
20'b01100100100101010010: color_data = 12'b000011110000;
20'b01100100100101010011: color_data = 12'b000011110000;
20'b01100100100101010100: color_data = 12'b000011110000;
20'b01100100100101010101: color_data = 12'b000011110000;
20'b01100100100101010110: color_data = 12'b000011110000;
20'b01100100100101010111: color_data = 12'b000011110000;
20'b01100100100101011000: color_data = 12'b000011110000;
20'b01100100100101011001: color_data = 12'b000011110000;
20'b01100100100101011010: color_data = 12'b000011110000;
20'b01100100100101011011: color_data = 12'b000011110000;
20'b01100100100101011100: color_data = 12'b000011110000;
20'b01100100100101011101: color_data = 12'b000011110000;
20'b01100100100101011110: color_data = 12'b000011110000;
20'b01100100100101011111: color_data = 12'b000011110000;
20'b01100100100101100011: color_data = 12'b111100001111;
20'b01100100100101100100: color_data = 12'b111100001111;
20'b01100100100101100101: color_data = 12'b111100001111;
20'b01100100100101100110: color_data = 12'b111100001111;
20'b01100100100101100111: color_data = 12'b111100001111;
20'b01100100100101101000: color_data = 12'b111100001111;
20'b01100100100101101001: color_data = 12'b111100001111;
20'b01100100100101101010: color_data = 12'b111100001111;
20'b01100100100101101011: color_data = 12'b111100001111;
20'b01100100100101101100: color_data = 12'b111100001111;
20'b01100100100101101101: color_data = 12'b111100001111;
20'b01100100100101101110: color_data = 12'b111100001111;
20'b01100100100101101111: color_data = 12'b111100001111;
20'b01100100100101110000: color_data = 12'b111100001111;
20'b01100100100101110001: color_data = 12'b111100001111;
20'b01100100100101110010: color_data = 12'b111100001111;
20'b01100100100101110011: color_data = 12'b111100001111;
20'b01100100100101110100: color_data = 12'b111100001111;
20'b01100100100101111000: color_data = 12'b111100001111;
20'b01100100100101111001: color_data = 12'b111100001111;
20'b01100100100101111010: color_data = 12'b111100001111;
20'b01100100100101111011: color_data = 12'b111100001111;
20'b01100100100101111100: color_data = 12'b111100001111;
20'b01100100100101111101: color_data = 12'b111100001111;
20'b01100100100101111110: color_data = 12'b111100001111;
20'b01100100100101111111: color_data = 12'b111100001111;
20'b01100100100110000000: color_data = 12'b111100001111;
20'b01100100100110000001: color_data = 12'b111100001111;
20'b01100100100110000010: color_data = 12'b111100001111;
20'b01100100100110000011: color_data = 12'b111100001111;
20'b01100100100110000100: color_data = 12'b111100001111;
20'b01100100100110000101: color_data = 12'b111100001111;
20'b01100100100110000110: color_data = 12'b111100001111;
20'b01100100100110000111: color_data = 12'b111100001111;
20'b01100100100110001000: color_data = 12'b111100001111;
20'b01100100100110001001: color_data = 12'b111100001111;
20'b01100100100110001101: color_data = 12'b111100000000;
20'b01100100100110001110: color_data = 12'b111100000000;
20'b01100100100110001111: color_data = 12'b111100000000;
20'b01100100100110010000: color_data = 12'b111100000000;
20'b01100100100110010001: color_data = 12'b111100000000;
20'b01100100100110010010: color_data = 12'b111100000000;
20'b01100100100110010011: color_data = 12'b111100000000;
20'b01100100100110010100: color_data = 12'b111100000000;
20'b01100100100110010101: color_data = 12'b111100000000;
20'b01100100100110010110: color_data = 12'b111100000000;
20'b01100100100110010111: color_data = 12'b111100000000;
20'b01100100100110011000: color_data = 12'b111100000000;
20'b01100100100110011001: color_data = 12'b111100000000;
20'b01100100100110011010: color_data = 12'b111100000000;
20'b01100100100110011011: color_data = 12'b111100000000;
20'b01100100100110011100: color_data = 12'b111100000000;
20'b01100100100110011101: color_data = 12'b111100000000;
20'b01100100100110011110: color_data = 12'b111100000000;
20'b01100100110011111010: color_data = 12'b000001101111;
20'b01100100110011111011: color_data = 12'b000001101111;
20'b01100100110011111100: color_data = 12'b000001101111;
20'b01100100110011111101: color_data = 12'b000001101111;
20'b01100100110011111110: color_data = 12'b000001101111;
20'b01100100110011111111: color_data = 12'b000001101111;
20'b01100100110100000000: color_data = 12'b000001101111;
20'b01100100110100000001: color_data = 12'b000001101111;
20'b01100100110100000010: color_data = 12'b000001101111;
20'b01100100110100000011: color_data = 12'b000001101111;
20'b01100100110100000100: color_data = 12'b000001101111;
20'b01100100110100000101: color_data = 12'b000001101111;
20'b01100100110100000110: color_data = 12'b000001101111;
20'b01100100110100000111: color_data = 12'b000001101111;
20'b01100100110100001000: color_data = 12'b000001101111;
20'b01100100110100001001: color_data = 12'b000001101111;
20'b01100100110100001010: color_data = 12'b000001101111;
20'b01100100110100001011: color_data = 12'b000001101111;
20'b01100100110100001111: color_data = 12'b000001101111;
20'b01100100110100010000: color_data = 12'b000001101111;
20'b01100100110100010001: color_data = 12'b000001101111;
20'b01100100110100010010: color_data = 12'b000001101111;
20'b01100100110100010011: color_data = 12'b000001101111;
20'b01100100110100010100: color_data = 12'b000001101111;
20'b01100100110100010101: color_data = 12'b000001101111;
20'b01100100110100010110: color_data = 12'b000001101111;
20'b01100100110100010111: color_data = 12'b000001101111;
20'b01100100110100011000: color_data = 12'b000001101111;
20'b01100100110100011001: color_data = 12'b000001101111;
20'b01100100110100011010: color_data = 12'b000001101111;
20'b01100100110100011011: color_data = 12'b000001101111;
20'b01100100110100011100: color_data = 12'b000001101111;
20'b01100100110100011101: color_data = 12'b000001101111;
20'b01100100110100011110: color_data = 12'b000001101111;
20'b01100100110100011111: color_data = 12'b000001101111;
20'b01100100110100100000: color_data = 12'b000001101111;
20'b01100100110100100100: color_data = 12'b000001101111;
20'b01100100110100100101: color_data = 12'b000001101111;
20'b01100100110100100110: color_data = 12'b000001101111;
20'b01100100110100100111: color_data = 12'b000001101111;
20'b01100100110100101000: color_data = 12'b000001101111;
20'b01100100110100101001: color_data = 12'b000001101111;
20'b01100100110100101010: color_data = 12'b000001101111;
20'b01100100110100101011: color_data = 12'b000001101111;
20'b01100100110100101100: color_data = 12'b000001101111;
20'b01100100110100101101: color_data = 12'b000001101111;
20'b01100100110100101110: color_data = 12'b000001101111;
20'b01100100110100101111: color_data = 12'b000001101111;
20'b01100100110100110000: color_data = 12'b000001101111;
20'b01100100110100110001: color_data = 12'b000001101111;
20'b01100100110100110010: color_data = 12'b000001101111;
20'b01100100110100110011: color_data = 12'b000001101111;
20'b01100100110100110100: color_data = 12'b000001101111;
20'b01100100110100110101: color_data = 12'b000001101111;
20'b01100100110100111001: color_data = 12'b000011110000;
20'b01100100110100111010: color_data = 12'b000011110000;
20'b01100100110100111011: color_data = 12'b000011110000;
20'b01100100110100111100: color_data = 12'b000011110000;
20'b01100100110100111101: color_data = 12'b000011110000;
20'b01100100110100111110: color_data = 12'b000011110000;
20'b01100100110100111111: color_data = 12'b000011110000;
20'b01100100110101000000: color_data = 12'b000011110000;
20'b01100100110101000001: color_data = 12'b000011110000;
20'b01100100110101000010: color_data = 12'b000011110000;
20'b01100100110101000011: color_data = 12'b000011110000;
20'b01100100110101000100: color_data = 12'b000011110000;
20'b01100100110101000101: color_data = 12'b000011110000;
20'b01100100110101000110: color_data = 12'b000011110000;
20'b01100100110101000111: color_data = 12'b000011110000;
20'b01100100110101001000: color_data = 12'b000011110000;
20'b01100100110101001001: color_data = 12'b000011110000;
20'b01100100110101001010: color_data = 12'b000011110000;
20'b01100100110101001110: color_data = 12'b000011110000;
20'b01100100110101001111: color_data = 12'b000011110000;
20'b01100100110101010000: color_data = 12'b000011110000;
20'b01100100110101010001: color_data = 12'b000011110000;
20'b01100100110101010010: color_data = 12'b000011110000;
20'b01100100110101010011: color_data = 12'b000011110000;
20'b01100100110101010100: color_data = 12'b000011110000;
20'b01100100110101010101: color_data = 12'b000011110000;
20'b01100100110101010110: color_data = 12'b000011110000;
20'b01100100110101010111: color_data = 12'b000011110000;
20'b01100100110101011000: color_data = 12'b000011110000;
20'b01100100110101011001: color_data = 12'b000011110000;
20'b01100100110101011010: color_data = 12'b000011110000;
20'b01100100110101011011: color_data = 12'b000011110000;
20'b01100100110101011100: color_data = 12'b000011110000;
20'b01100100110101011101: color_data = 12'b000011110000;
20'b01100100110101011110: color_data = 12'b000011110000;
20'b01100100110101011111: color_data = 12'b000011110000;
20'b01100100110101100011: color_data = 12'b111100001111;
20'b01100100110101100100: color_data = 12'b111100001111;
20'b01100100110101100101: color_data = 12'b111100001111;
20'b01100100110101100110: color_data = 12'b111100001111;
20'b01100100110101100111: color_data = 12'b111100001111;
20'b01100100110101101000: color_data = 12'b111100001111;
20'b01100100110101101001: color_data = 12'b111100001111;
20'b01100100110101101010: color_data = 12'b111100001111;
20'b01100100110101101011: color_data = 12'b111100001111;
20'b01100100110101101100: color_data = 12'b111100001111;
20'b01100100110101101101: color_data = 12'b111100001111;
20'b01100100110101101110: color_data = 12'b111100001111;
20'b01100100110101101111: color_data = 12'b111100001111;
20'b01100100110101110000: color_data = 12'b111100001111;
20'b01100100110101110001: color_data = 12'b111100001111;
20'b01100100110101110010: color_data = 12'b111100001111;
20'b01100100110101110011: color_data = 12'b111100001111;
20'b01100100110101110100: color_data = 12'b111100001111;
20'b01100100110101111000: color_data = 12'b111100001111;
20'b01100100110101111001: color_data = 12'b111100001111;
20'b01100100110101111010: color_data = 12'b111100001111;
20'b01100100110101111011: color_data = 12'b111100001111;
20'b01100100110101111100: color_data = 12'b111100001111;
20'b01100100110101111101: color_data = 12'b111100001111;
20'b01100100110101111110: color_data = 12'b111100001111;
20'b01100100110101111111: color_data = 12'b111100001111;
20'b01100100110110000000: color_data = 12'b111100001111;
20'b01100100110110000001: color_data = 12'b111100001111;
20'b01100100110110000010: color_data = 12'b111100001111;
20'b01100100110110000011: color_data = 12'b111100001111;
20'b01100100110110000100: color_data = 12'b111100001111;
20'b01100100110110000101: color_data = 12'b111100001111;
20'b01100100110110000110: color_data = 12'b111100001111;
20'b01100100110110000111: color_data = 12'b111100001111;
20'b01100100110110001000: color_data = 12'b111100001111;
20'b01100100110110001001: color_data = 12'b111100001111;
20'b01100100110110001101: color_data = 12'b111100000000;
20'b01100100110110001110: color_data = 12'b111100000000;
20'b01100100110110001111: color_data = 12'b111100000000;
20'b01100100110110010000: color_data = 12'b111100000000;
20'b01100100110110010001: color_data = 12'b111100000000;
20'b01100100110110010010: color_data = 12'b111100000000;
20'b01100100110110010011: color_data = 12'b111100000000;
20'b01100100110110010100: color_data = 12'b111100000000;
20'b01100100110110010101: color_data = 12'b111100000000;
20'b01100100110110010110: color_data = 12'b111100000000;
20'b01100100110110010111: color_data = 12'b111100000000;
20'b01100100110110011000: color_data = 12'b111100000000;
20'b01100100110110011001: color_data = 12'b111100000000;
20'b01100100110110011010: color_data = 12'b111100000000;
20'b01100100110110011011: color_data = 12'b111100000000;
20'b01100100110110011100: color_data = 12'b111100000000;
20'b01100100110110011101: color_data = 12'b111100000000;
20'b01100100110110011110: color_data = 12'b111100000000;
20'b01100101000011111010: color_data = 12'b000001101111;
20'b01100101000011111011: color_data = 12'b000001101111;
20'b01100101000011111100: color_data = 12'b000001101111;
20'b01100101000011111101: color_data = 12'b000001101111;
20'b01100101000011111110: color_data = 12'b000001101111;
20'b01100101000011111111: color_data = 12'b000001101111;
20'b01100101000100000000: color_data = 12'b000001101111;
20'b01100101000100000001: color_data = 12'b000001101111;
20'b01100101000100000010: color_data = 12'b000001101111;
20'b01100101000100000011: color_data = 12'b000001101111;
20'b01100101000100000100: color_data = 12'b000001101111;
20'b01100101000100000101: color_data = 12'b000001101111;
20'b01100101000100000110: color_data = 12'b000001101111;
20'b01100101000100000111: color_data = 12'b000001101111;
20'b01100101000100001000: color_data = 12'b000001101111;
20'b01100101000100001001: color_data = 12'b000001101111;
20'b01100101000100001010: color_data = 12'b000001101111;
20'b01100101000100001011: color_data = 12'b000001101111;
20'b01100101000100001111: color_data = 12'b000001101111;
20'b01100101000100010000: color_data = 12'b000001101111;
20'b01100101000100010001: color_data = 12'b000001101111;
20'b01100101000100010010: color_data = 12'b000001101111;
20'b01100101000100010011: color_data = 12'b000001101111;
20'b01100101000100010100: color_data = 12'b000001101111;
20'b01100101000100010101: color_data = 12'b000001101111;
20'b01100101000100010110: color_data = 12'b000001101111;
20'b01100101000100010111: color_data = 12'b000001101111;
20'b01100101000100011000: color_data = 12'b000001101111;
20'b01100101000100011001: color_data = 12'b000001101111;
20'b01100101000100011010: color_data = 12'b000001101111;
20'b01100101000100011011: color_data = 12'b000001101111;
20'b01100101000100011100: color_data = 12'b000001101111;
20'b01100101000100011101: color_data = 12'b000001101111;
20'b01100101000100011110: color_data = 12'b000001101111;
20'b01100101000100011111: color_data = 12'b000001101111;
20'b01100101000100100000: color_data = 12'b000001101111;
20'b01100101000100100100: color_data = 12'b000001101111;
20'b01100101000100100101: color_data = 12'b000001101111;
20'b01100101000100100110: color_data = 12'b000001101111;
20'b01100101000100100111: color_data = 12'b000001101111;
20'b01100101000100101000: color_data = 12'b000001101111;
20'b01100101000100101001: color_data = 12'b000001101111;
20'b01100101000100101010: color_data = 12'b000001101111;
20'b01100101000100101011: color_data = 12'b000001101111;
20'b01100101000100101100: color_data = 12'b000001101111;
20'b01100101000100101101: color_data = 12'b000001101111;
20'b01100101000100101110: color_data = 12'b000001101111;
20'b01100101000100101111: color_data = 12'b000001101111;
20'b01100101000100110000: color_data = 12'b000001101111;
20'b01100101000100110001: color_data = 12'b000001101111;
20'b01100101000100110010: color_data = 12'b000001101111;
20'b01100101000100110011: color_data = 12'b000001101111;
20'b01100101000100110100: color_data = 12'b000001101111;
20'b01100101000100110101: color_data = 12'b000001101111;
20'b01100101000100111001: color_data = 12'b000011110000;
20'b01100101000100111010: color_data = 12'b000011110000;
20'b01100101000100111011: color_data = 12'b000011110000;
20'b01100101000100111100: color_data = 12'b000011110000;
20'b01100101000100111101: color_data = 12'b000011110000;
20'b01100101000100111110: color_data = 12'b000011110000;
20'b01100101000100111111: color_data = 12'b000011110000;
20'b01100101000101000000: color_data = 12'b000011110000;
20'b01100101000101000001: color_data = 12'b000011110000;
20'b01100101000101000010: color_data = 12'b000011110000;
20'b01100101000101000011: color_data = 12'b000011110000;
20'b01100101000101000100: color_data = 12'b000011110000;
20'b01100101000101000101: color_data = 12'b000011110000;
20'b01100101000101000110: color_data = 12'b000011110000;
20'b01100101000101000111: color_data = 12'b000011110000;
20'b01100101000101001000: color_data = 12'b000011110000;
20'b01100101000101001001: color_data = 12'b000011110000;
20'b01100101000101001010: color_data = 12'b000011110000;
20'b01100101000101001110: color_data = 12'b000011110000;
20'b01100101000101001111: color_data = 12'b000011110000;
20'b01100101000101010000: color_data = 12'b000011110000;
20'b01100101000101010001: color_data = 12'b000011110000;
20'b01100101000101010010: color_data = 12'b000011110000;
20'b01100101000101010011: color_data = 12'b000011110000;
20'b01100101000101010100: color_data = 12'b000011110000;
20'b01100101000101010101: color_data = 12'b000011110000;
20'b01100101000101010110: color_data = 12'b000011110000;
20'b01100101000101010111: color_data = 12'b000011110000;
20'b01100101000101011000: color_data = 12'b000011110000;
20'b01100101000101011001: color_data = 12'b000011110000;
20'b01100101000101011010: color_data = 12'b000011110000;
20'b01100101000101011011: color_data = 12'b000011110000;
20'b01100101000101011100: color_data = 12'b000011110000;
20'b01100101000101011101: color_data = 12'b000011110000;
20'b01100101000101011110: color_data = 12'b000011110000;
20'b01100101000101011111: color_data = 12'b000011110000;
20'b01100101000101100011: color_data = 12'b111100001111;
20'b01100101000101100100: color_data = 12'b111100001111;
20'b01100101000101100101: color_data = 12'b111100001111;
20'b01100101000101100110: color_data = 12'b111100001111;
20'b01100101000101100111: color_data = 12'b111100001111;
20'b01100101000101101000: color_data = 12'b111100001111;
20'b01100101000101101001: color_data = 12'b111100001111;
20'b01100101000101101010: color_data = 12'b111100001111;
20'b01100101000101101011: color_data = 12'b111100001111;
20'b01100101000101101100: color_data = 12'b111100001111;
20'b01100101000101101101: color_data = 12'b111100001111;
20'b01100101000101101110: color_data = 12'b111100001111;
20'b01100101000101101111: color_data = 12'b111100001111;
20'b01100101000101110000: color_data = 12'b111100001111;
20'b01100101000101110001: color_data = 12'b111100001111;
20'b01100101000101110010: color_data = 12'b111100001111;
20'b01100101000101110011: color_data = 12'b111100001111;
20'b01100101000101110100: color_data = 12'b111100001111;
20'b01100101000101111000: color_data = 12'b111100001111;
20'b01100101000101111001: color_data = 12'b111100001111;
20'b01100101000101111010: color_data = 12'b111100001111;
20'b01100101000101111011: color_data = 12'b111100001111;
20'b01100101000101111100: color_data = 12'b111100001111;
20'b01100101000101111101: color_data = 12'b111100001111;
20'b01100101000101111110: color_data = 12'b111100001111;
20'b01100101000101111111: color_data = 12'b111100001111;
20'b01100101000110000000: color_data = 12'b111100001111;
20'b01100101000110000001: color_data = 12'b111100001111;
20'b01100101000110000010: color_data = 12'b111100001111;
20'b01100101000110000011: color_data = 12'b111100001111;
20'b01100101000110000100: color_data = 12'b111100001111;
20'b01100101000110000101: color_data = 12'b111100001111;
20'b01100101000110000110: color_data = 12'b111100001111;
20'b01100101000110000111: color_data = 12'b111100001111;
20'b01100101000110001000: color_data = 12'b111100001111;
20'b01100101000110001001: color_data = 12'b111100001111;
20'b01100101000110001101: color_data = 12'b111100000000;
20'b01100101000110001110: color_data = 12'b111100000000;
20'b01100101000110001111: color_data = 12'b111100000000;
20'b01100101000110010000: color_data = 12'b111100000000;
20'b01100101000110010001: color_data = 12'b111100000000;
20'b01100101000110010010: color_data = 12'b111100000000;
20'b01100101000110010011: color_data = 12'b111100000000;
20'b01100101000110010100: color_data = 12'b111100000000;
20'b01100101000110010101: color_data = 12'b111100000000;
20'b01100101000110010110: color_data = 12'b111100000000;
20'b01100101000110010111: color_data = 12'b111100000000;
20'b01100101000110011000: color_data = 12'b111100000000;
20'b01100101000110011001: color_data = 12'b111100000000;
20'b01100101000110011010: color_data = 12'b111100000000;
20'b01100101000110011011: color_data = 12'b111100000000;
20'b01100101000110011100: color_data = 12'b111100000000;
20'b01100101000110011101: color_data = 12'b111100000000;
20'b01100101000110011110: color_data = 12'b111100000000;
20'b01100101010011111010: color_data = 12'b000001101111;
20'b01100101010011111011: color_data = 12'b000001101111;
20'b01100101010011111100: color_data = 12'b000001101111;
20'b01100101010011111101: color_data = 12'b000001101111;
20'b01100101010011111110: color_data = 12'b000001101111;
20'b01100101010011111111: color_data = 12'b000001101111;
20'b01100101010100000000: color_data = 12'b000001101111;
20'b01100101010100000001: color_data = 12'b000001101111;
20'b01100101010100000010: color_data = 12'b000001101111;
20'b01100101010100000011: color_data = 12'b000001101111;
20'b01100101010100000100: color_data = 12'b000001101111;
20'b01100101010100000101: color_data = 12'b000001101111;
20'b01100101010100000110: color_data = 12'b000001101111;
20'b01100101010100000111: color_data = 12'b000001101111;
20'b01100101010100001000: color_data = 12'b000001101111;
20'b01100101010100001001: color_data = 12'b000001101111;
20'b01100101010100001010: color_data = 12'b000001101111;
20'b01100101010100001011: color_data = 12'b000001101111;
20'b01100101010100001111: color_data = 12'b000001101111;
20'b01100101010100010000: color_data = 12'b000001101111;
20'b01100101010100010001: color_data = 12'b000001101111;
20'b01100101010100010010: color_data = 12'b000001101111;
20'b01100101010100010011: color_data = 12'b000001101111;
20'b01100101010100010100: color_data = 12'b000001101111;
20'b01100101010100010101: color_data = 12'b000001101111;
20'b01100101010100010110: color_data = 12'b000001101111;
20'b01100101010100010111: color_data = 12'b000001101111;
20'b01100101010100011000: color_data = 12'b000001101111;
20'b01100101010100011001: color_data = 12'b000001101111;
20'b01100101010100011010: color_data = 12'b000001101111;
20'b01100101010100011011: color_data = 12'b000001101111;
20'b01100101010100011100: color_data = 12'b000001101111;
20'b01100101010100011101: color_data = 12'b000001101111;
20'b01100101010100011110: color_data = 12'b000001101111;
20'b01100101010100011111: color_data = 12'b000001101111;
20'b01100101010100100000: color_data = 12'b000001101111;
20'b01100101010100100100: color_data = 12'b000001101111;
20'b01100101010100100101: color_data = 12'b000001101111;
20'b01100101010100100110: color_data = 12'b000001101111;
20'b01100101010100100111: color_data = 12'b000001101111;
20'b01100101010100101000: color_data = 12'b000001101111;
20'b01100101010100101001: color_data = 12'b000001101111;
20'b01100101010100101010: color_data = 12'b000001101111;
20'b01100101010100101011: color_data = 12'b000001101111;
20'b01100101010100101100: color_data = 12'b000001101111;
20'b01100101010100101101: color_data = 12'b000001101111;
20'b01100101010100101110: color_data = 12'b000001101111;
20'b01100101010100101111: color_data = 12'b000001101111;
20'b01100101010100110000: color_data = 12'b000001101111;
20'b01100101010100110001: color_data = 12'b000001101111;
20'b01100101010100110010: color_data = 12'b000001101111;
20'b01100101010100110011: color_data = 12'b000001101111;
20'b01100101010100110100: color_data = 12'b000001101111;
20'b01100101010100110101: color_data = 12'b000001101111;
20'b01100101010100111001: color_data = 12'b000011110000;
20'b01100101010100111010: color_data = 12'b000011110000;
20'b01100101010100111011: color_data = 12'b000011110000;
20'b01100101010100111100: color_data = 12'b000011110000;
20'b01100101010100111101: color_data = 12'b000011110000;
20'b01100101010100111110: color_data = 12'b000011110000;
20'b01100101010100111111: color_data = 12'b000011110000;
20'b01100101010101000000: color_data = 12'b000011110000;
20'b01100101010101000001: color_data = 12'b000011110000;
20'b01100101010101000010: color_data = 12'b000011110000;
20'b01100101010101000011: color_data = 12'b000011110000;
20'b01100101010101000100: color_data = 12'b000011110000;
20'b01100101010101000101: color_data = 12'b000011110000;
20'b01100101010101000110: color_data = 12'b000011110000;
20'b01100101010101000111: color_data = 12'b000011110000;
20'b01100101010101001000: color_data = 12'b000011110000;
20'b01100101010101001001: color_data = 12'b000011110000;
20'b01100101010101001010: color_data = 12'b000011110000;
20'b01100101010101001110: color_data = 12'b000011110000;
20'b01100101010101001111: color_data = 12'b000011110000;
20'b01100101010101010000: color_data = 12'b000011110000;
20'b01100101010101010001: color_data = 12'b000011110000;
20'b01100101010101010010: color_data = 12'b000011110000;
20'b01100101010101010011: color_data = 12'b000011110000;
20'b01100101010101010100: color_data = 12'b000011110000;
20'b01100101010101010101: color_data = 12'b000011110000;
20'b01100101010101010110: color_data = 12'b000011110000;
20'b01100101010101010111: color_data = 12'b000011110000;
20'b01100101010101011000: color_data = 12'b000011110000;
20'b01100101010101011001: color_data = 12'b000011110000;
20'b01100101010101011010: color_data = 12'b000011110000;
20'b01100101010101011011: color_data = 12'b000011110000;
20'b01100101010101011100: color_data = 12'b000011110000;
20'b01100101010101011101: color_data = 12'b000011110000;
20'b01100101010101011110: color_data = 12'b000011110000;
20'b01100101010101011111: color_data = 12'b000011110000;
20'b01100101010101100011: color_data = 12'b111100001111;
20'b01100101010101100100: color_data = 12'b111100001111;
20'b01100101010101100101: color_data = 12'b111100001111;
20'b01100101010101100110: color_data = 12'b111100001111;
20'b01100101010101100111: color_data = 12'b111100001111;
20'b01100101010101101000: color_data = 12'b111100001111;
20'b01100101010101101001: color_data = 12'b111100001111;
20'b01100101010101101010: color_data = 12'b111100001111;
20'b01100101010101101011: color_data = 12'b111100001111;
20'b01100101010101101100: color_data = 12'b111100001111;
20'b01100101010101101101: color_data = 12'b111100001111;
20'b01100101010101101110: color_data = 12'b111100001111;
20'b01100101010101101111: color_data = 12'b111100001111;
20'b01100101010101110000: color_data = 12'b111100001111;
20'b01100101010101110001: color_data = 12'b111100001111;
20'b01100101010101110010: color_data = 12'b111100001111;
20'b01100101010101110011: color_data = 12'b111100001111;
20'b01100101010101110100: color_data = 12'b111100001111;
20'b01100101010101111000: color_data = 12'b111100001111;
20'b01100101010101111001: color_data = 12'b111100001111;
20'b01100101010101111010: color_data = 12'b111100001111;
20'b01100101010101111011: color_data = 12'b111100001111;
20'b01100101010101111100: color_data = 12'b111100001111;
20'b01100101010101111101: color_data = 12'b111100001111;
20'b01100101010101111110: color_data = 12'b111100001111;
20'b01100101010101111111: color_data = 12'b111100001111;
20'b01100101010110000000: color_data = 12'b111100001111;
20'b01100101010110000001: color_data = 12'b111100001111;
20'b01100101010110000010: color_data = 12'b111100001111;
20'b01100101010110000011: color_data = 12'b111100001111;
20'b01100101010110000100: color_data = 12'b111100001111;
20'b01100101010110000101: color_data = 12'b111100001111;
20'b01100101010110000110: color_data = 12'b111100001111;
20'b01100101010110000111: color_data = 12'b111100001111;
20'b01100101010110001000: color_data = 12'b111100001111;
20'b01100101010110001001: color_data = 12'b111100001111;
20'b01100101010110001101: color_data = 12'b111100000000;
20'b01100101010110001110: color_data = 12'b111100000000;
20'b01100101010110001111: color_data = 12'b111100000000;
20'b01100101010110010000: color_data = 12'b111100000000;
20'b01100101010110010001: color_data = 12'b111100000000;
20'b01100101010110010010: color_data = 12'b111100000000;
20'b01100101010110010011: color_data = 12'b111100000000;
20'b01100101010110010100: color_data = 12'b111100000000;
20'b01100101010110010101: color_data = 12'b111100000000;
20'b01100101010110010110: color_data = 12'b111100000000;
20'b01100101010110010111: color_data = 12'b111100000000;
20'b01100101010110011000: color_data = 12'b111100000000;
20'b01100101010110011001: color_data = 12'b111100000000;
20'b01100101010110011010: color_data = 12'b111100000000;
20'b01100101010110011011: color_data = 12'b111100000000;
20'b01100101010110011100: color_data = 12'b111100000000;
20'b01100101010110011101: color_data = 12'b111100000000;
20'b01100101010110011110: color_data = 12'b111100000000;
20'b01100101100011111010: color_data = 12'b000001101111;
20'b01100101100011111011: color_data = 12'b000001101111;
20'b01100101100011111100: color_data = 12'b000001101111;
20'b01100101100011111101: color_data = 12'b000001101111;
20'b01100101100011111110: color_data = 12'b000001101111;
20'b01100101100011111111: color_data = 12'b000001101111;
20'b01100101100100000000: color_data = 12'b000001101111;
20'b01100101100100000001: color_data = 12'b000001101111;
20'b01100101100100000010: color_data = 12'b000001101111;
20'b01100101100100000011: color_data = 12'b000001101111;
20'b01100101100100000100: color_data = 12'b000001101111;
20'b01100101100100000101: color_data = 12'b000001101111;
20'b01100101100100000110: color_data = 12'b000001101111;
20'b01100101100100000111: color_data = 12'b000001101111;
20'b01100101100100001000: color_data = 12'b000001101111;
20'b01100101100100001001: color_data = 12'b000001101111;
20'b01100101100100001010: color_data = 12'b000001101111;
20'b01100101100100001011: color_data = 12'b000001101111;
20'b01100101100100001111: color_data = 12'b000001101111;
20'b01100101100100010000: color_data = 12'b000001101111;
20'b01100101100100010001: color_data = 12'b000001101111;
20'b01100101100100010010: color_data = 12'b000001101111;
20'b01100101100100010011: color_data = 12'b000001101111;
20'b01100101100100010100: color_data = 12'b000001101111;
20'b01100101100100010101: color_data = 12'b000001101111;
20'b01100101100100010110: color_data = 12'b000001101111;
20'b01100101100100010111: color_data = 12'b000001101111;
20'b01100101100100011000: color_data = 12'b000001101111;
20'b01100101100100011001: color_data = 12'b000001101111;
20'b01100101100100011010: color_data = 12'b000001101111;
20'b01100101100100011011: color_data = 12'b000001101111;
20'b01100101100100011100: color_data = 12'b000001101111;
20'b01100101100100011101: color_data = 12'b000001101111;
20'b01100101100100011110: color_data = 12'b000001101111;
20'b01100101100100011111: color_data = 12'b000001101111;
20'b01100101100100100000: color_data = 12'b000001101111;
20'b01100101100100100100: color_data = 12'b000001101111;
20'b01100101100100100101: color_data = 12'b000001101111;
20'b01100101100100100110: color_data = 12'b000001101111;
20'b01100101100100100111: color_data = 12'b000001101111;
20'b01100101100100101000: color_data = 12'b000001101111;
20'b01100101100100101001: color_data = 12'b000001101111;
20'b01100101100100101010: color_data = 12'b000001101111;
20'b01100101100100101011: color_data = 12'b000001101111;
20'b01100101100100101100: color_data = 12'b000001101111;
20'b01100101100100101101: color_data = 12'b000001101111;
20'b01100101100100101110: color_data = 12'b000001101111;
20'b01100101100100101111: color_data = 12'b000001101111;
20'b01100101100100110000: color_data = 12'b000001101111;
20'b01100101100100110001: color_data = 12'b000001101111;
20'b01100101100100110010: color_data = 12'b000001101111;
20'b01100101100100110011: color_data = 12'b000001101111;
20'b01100101100100110100: color_data = 12'b000001101111;
20'b01100101100100110101: color_data = 12'b000001101111;
20'b01100101100100111001: color_data = 12'b000011110000;
20'b01100101100100111010: color_data = 12'b000011110000;
20'b01100101100100111011: color_data = 12'b000011110000;
20'b01100101100100111100: color_data = 12'b000011110000;
20'b01100101100100111101: color_data = 12'b000011110000;
20'b01100101100100111110: color_data = 12'b000011110000;
20'b01100101100100111111: color_data = 12'b000011110000;
20'b01100101100101000000: color_data = 12'b000011110000;
20'b01100101100101000001: color_data = 12'b000011110000;
20'b01100101100101000010: color_data = 12'b000011110000;
20'b01100101100101000011: color_data = 12'b000011110000;
20'b01100101100101000100: color_data = 12'b000011110000;
20'b01100101100101000101: color_data = 12'b000011110000;
20'b01100101100101000110: color_data = 12'b000011110000;
20'b01100101100101000111: color_data = 12'b000011110000;
20'b01100101100101001000: color_data = 12'b000011110000;
20'b01100101100101001001: color_data = 12'b000011110000;
20'b01100101100101001010: color_data = 12'b000011110000;
20'b01100101100101001110: color_data = 12'b000011110000;
20'b01100101100101001111: color_data = 12'b000011110000;
20'b01100101100101010000: color_data = 12'b000011110000;
20'b01100101100101010001: color_data = 12'b000011110000;
20'b01100101100101010010: color_data = 12'b000011110000;
20'b01100101100101010011: color_data = 12'b000011110000;
20'b01100101100101010100: color_data = 12'b000011110000;
20'b01100101100101010101: color_data = 12'b000011110000;
20'b01100101100101010110: color_data = 12'b000011110000;
20'b01100101100101010111: color_data = 12'b000011110000;
20'b01100101100101011000: color_data = 12'b000011110000;
20'b01100101100101011001: color_data = 12'b000011110000;
20'b01100101100101011010: color_data = 12'b000011110000;
20'b01100101100101011011: color_data = 12'b000011110000;
20'b01100101100101011100: color_data = 12'b000011110000;
20'b01100101100101011101: color_data = 12'b000011110000;
20'b01100101100101011110: color_data = 12'b000011110000;
20'b01100101100101011111: color_data = 12'b000011110000;
20'b01100101100101100011: color_data = 12'b111100001111;
20'b01100101100101100100: color_data = 12'b111100001111;
20'b01100101100101100101: color_data = 12'b111100001111;
20'b01100101100101100110: color_data = 12'b111100001111;
20'b01100101100101100111: color_data = 12'b111100001111;
20'b01100101100101101000: color_data = 12'b111100001111;
20'b01100101100101101001: color_data = 12'b111100001111;
20'b01100101100101101010: color_data = 12'b111100001111;
20'b01100101100101101011: color_data = 12'b111100001111;
20'b01100101100101101100: color_data = 12'b111100001111;
20'b01100101100101101101: color_data = 12'b111100001111;
20'b01100101100101101110: color_data = 12'b111100001111;
20'b01100101100101101111: color_data = 12'b111100001111;
20'b01100101100101110000: color_data = 12'b111100001111;
20'b01100101100101110001: color_data = 12'b111100001111;
20'b01100101100101110010: color_data = 12'b111100001111;
20'b01100101100101110011: color_data = 12'b111100001111;
20'b01100101100101110100: color_data = 12'b111100001111;
20'b01100101100101111000: color_data = 12'b111100001111;
20'b01100101100101111001: color_data = 12'b111100001111;
20'b01100101100101111010: color_data = 12'b111100001111;
20'b01100101100101111011: color_data = 12'b111100001111;
20'b01100101100101111100: color_data = 12'b111100001111;
20'b01100101100101111101: color_data = 12'b111100001111;
20'b01100101100101111110: color_data = 12'b111100001111;
20'b01100101100101111111: color_data = 12'b111100001111;
20'b01100101100110000000: color_data = 12'b111100001111;
20'b01100101100110000001: color_data = 12'b111100001111;
20'b01100101100110000010: color_data = 12'b111100001111;
20'b01100101100110000011: color_data = 12'b111100001111;
20'b01100101100110000100: color_data = 12'b111100001111;
20'b01100101100110000101: color_data = 12'b111100001111;
20'b01100101100110000110: color_data = 12'b111100001111;
20'b01100101100110000111: color_data = 12'b111100001111;
20'b01100101100110001000: color_data = 12'b111100001111;
20'b01100101100110001001: color_data = 12'b111100001111;
20'b01100101100110001101: color_data = 12'b111100000000;
20'b01100101100110001110: color_data = 12'b111100000000;
20'b01100101100110001111: color_data = 12'b111100000000;
20'b01100101100110010000: color_data = 12'b111100000000;
20'b01100101100110010001: color_data = 12'b111100000000;
20'b01100101100110010010: color_data = 12'b111100000000;
20'b01100101100110010011: color_data = 12'b111100000000;
20'b01100101100110010100: color_data = 12'b111100000000;
20'b01100101100110010101: color_data = 12'b111100000000;
20'b01100101100110010110: color_data = 12'b111100000000;
20'b01100101100110010111: color_data = 12'b111100000000;
20'b01100101100110011000: color_data = 12'b111100000000;
20'b01100101100110011001: color_data = 12'b111100000000;
20'b01100101100110011010: color_data = 12'b111100000000;
20'b01100101100110011011: color_data = 12'b111100000000;
20'b01100101100110011100: color_data = 12'b111100000000;
20'b01100101100110011101: color_data = 12'b111100000000;
20'b01100101100110011110: color_data = 12'b111100000000;
20'b01100101110011111010: color_data = 12'b000001101111;
20'b01100101110011111011: color_data = 12'b000001101111;
20'b01100101110011111100: color_data = 12'b000001101111;
20'b01100101110011111101: color_data = 12'b000001101111;
20'b01100101110011111110: color_data = 12'b000001101111;
20'b01100101110011111111: color_data = 12'b000001101111;
20'b01100101110100000000: color_data = 12'b000001101111;
20'b01100101110100000001: color_data = 12'b000001101111;
20'b01100101110100000010: color_data = 12'b000001101111;
20'b01100101110100000011: color_data = 12'b000001101111;
20'b01100101110100000100: color_data = 12'b000001101111;
20'b01100101110100000101: color_data = 12'b000001101111;
20'b01100101110100000110: color_data = 12'b000001101111;
20'b01100101110100000111: color_data = 12'b000001101111;
20'b01100101110100001000: color_data = 12'b000001101111;
20'b01100101110100001001: color_data = 12'b000001101111;
20'b01100101110100001010: color_data = 12'b000001101111;
20'b01100101110100001011: color_data = 12'b000001101111;
20'b01100101110100001111: color_data = 12'b000001101111;
20'b01100101110100010000: color_data = 12'b000001101111;
20'b01100101110100010001: color_data = 12'b000001101111;
20'b01100101110100010010: color_data = 12'b000001101111;
20'b01100101110100010011: color_data = 12'b000001101111;
20'b01100101110100010100: color_data = 12'b000001101111;
20'b01100101110100010101: color_data = 12'b000001101111;
20'b01100101110100010110: color_data = 12'b000001101111;
20'b01100101110100010111: color_data = 12'b000001101111;
20'b01100101110100011000: color_data = 12'b000001101111;
20'b01100101110100011001: color_data = 12'b000001101111;
20'b01100101110100011010: color_data = 12'b000001101111;
20'b01100101110100011011: color_data = 12'b000001101111;
20'b01100101110100011100: color_data = 12'b000001101111;
20'b01100101110100011101: color_data = 12'b000001101111;
20'b01100101110100011110: color_data = 12'b000001101111;
20'b01100101110100011111: color_data = 12'b000001101111;
20'b01100101110100100000: color_data = 12'b000001101111;
20'b01100101110100100100: color_data = 12'b000001101111;
20'b01100101110100100101: color_data = 12'b000001101111;
20'b01100101110100100110: color_data = 12'b000001101111;
20'b01100101110100100111: color_data = 12'b000001101111;
20'b01100101110100101000: color_data = 12'b000001101111;
20'b01100101110100101001: color_data = 12'b000001101111;
20'b01100101110100101010: color_data = 12'b000001101111;
20'b01100101110100101011: color_data = 12'b000001101111;
20'b01100101110100101100: color_data = 12'b000001101111;
20'b01100101110100101101: color_data = 12'b000001101111;
20'b01100101110100101110: color_data = 12'b000001101111;
20'b01100101110100101111: color_data = 12'b000001101111;
20'b01100101110100110000: color_data = 12'b000001101111;
20'b01100101110100110001: color_data = 12'b000001101111;
20'b01100101110100110010: color_data = 12'b000001101111;
20'b01100101110100110011: color_data = 12'b000001101111;
20'b01100101110100110100: color_data = 12'b000001101111;
20'b01100101110100110101: color_data = 12'b000001101111;
20'b01100101110100111001: color_data = 12'b000011110000;
20'b01100101110100111010: color_data = 12'b000011110000;
20'b01100101110100111011: color_data = 12'b000011110000;
20'b01100101110100111100: color_data = 12'b000011110000;
20'b01100101110100111101: color_data = 12'b000011110000;
20'b01100101110100111110: color_data = 12'b000011110000;
20'b01100101110100111111: color_data = 12'b000011110000;
20'b01100101110101000000: color_data = 12'b000011110000;
20'b01100101110101000001: color_data = 12'b000011110000;
20'b01100101110101000010: color_data = 12'b000011110000;
20'b01100101110101000011: color_data = 12'b000011110000;
20'b01100101110101000100: color_data = 12'b000011110000;
20'b01100101110101000101: color_data = 12'b000011110000;
20'b01100101110101000110: color_data = 12'b000011110000;
20'b01100101110101000111: color_data = 12'b000011110000;
20'b01100101110101001000: color_data = 12'b000011110000;
20'b01100101110101001001: color_data = 12'b000011110000;
20'b01100101110101001010: color_data = 12'b000011110000;
20'b01100101110101001110: color_data = 12'b000011110000;
20'b01100101110101001111: color_data = 12'b000011110000;
20'b01100101110101010000: color_data = 12'b000011110000;
20'b01100101110101010001: color_data = 12'b000011110000;
20'b01100101110101010010: color_data = 12'b000011110000;
20'b01100101110101010011: color_data = 12'b000011110000;
20'b01100101110101010100: color_data = 12'b000011110000;
20'b01100101110101010101: color_data = 12'b000011110000;
20'b01100101110101010110: color_data = 12'b000011110000;
20'b01100101110101010111: color_data = 12'b000011110000;
20'b01100101110101011000: color_data = 12'b000011110000;
20'b01100101110101011001: color_data = 12'b000011110000;
20'b01100101110101011010: color_data = 12'b000011110000;
20'b01100101110101011011: color_data = 12'b000011110000;
20'b01100101110101011100: color_data = 12'b000011110000;
20'b01100101110101011101: color_data = 12'b000011110000;
20'b01100101110101011110: color_data = 12'b000011110000;
20'b01100101110101011111: color_data = 12'b000011110000;
20'b01100101110101100011: color_data = 12'b111100001111;
20'b01100101110101100100: color_data = 12'b111100001111;
20'b01100101110101100101: color_data = 12'b111100001111;
20'b01100101110101100110: color_data = 12'b111100001111;
20'b01100101110101100111: color_data = 12'b111100001111;
20'b01100101110101101000: color_data = 12'b111100001111;
20'b01100101110101101001: color_data = 12'b111100001111;
20'b01100101110101101010: color_data = 12'b111100001111;
20'b01100101110101101011: color_data = 12'b111100001111;
20'b01100101110101101100: color_data = 12'b111100001111;
20'b01100101110101101101: color_data = 12'b111100001111;
20'b01100101110101101110: color_data = 12'b111100001111;
20'b01100101110101101111: color_data = 12'b111100001111;
20'b01100101110101110000: color_data = 12'b111100001111;
20'b01100101110101110001: color_data = 12'b111100001111;
20'b01100101110101110010: color_data = 12'b111100001111;
20'b01100101110101110011: color_data = 12'b111100001111;
20'b01100101110101110100: color_data = 12'b111100001111;
20'b01100101110101111000: color_data = 12'b111100001111;
20'b01100101110101111001: color_data = 12'b111100001111;
20'b01100101110101111010: color_data = 12'b111100001111;
20'b01100101110101111011: color_data = 12'b111100001111;
20'b01100101110101111100: color_data = 12'b111100001111;
20'b01100101110101111101: color_data = 12'b111100001111;
20'b01100101110101111110: color_data = 12'b111100001111;
20'b01100101110101111111: color_data = 12'b111100001111;
20'b01100101110110000000: color_data = 12'b111100001111;
20'b01100101110110000001: color_data = 12'b111100001111;
20'b01100101110110000010: color_data = 12'b111100001111;
20'b01100101110110000011: color_data = 12'b111100001111;
20'b01100101110110000100: color_data = 12'b111100001111;
20'b01100101110110000101: color_data = 12'b111100001111;
20'b01100101110110000110: color_data = 12'b111100001111;
20'b01100101110110000111: color_data = 12'b111100001111;
20'b01100101110110001000: color_data = 12'b111100001111;
20'b01100101110110001001: color_data = 12'b111100001111;
20'b01100101110110001101: color_data = 12'b111100000000;
20'b01100101110110001110: color_data = 12'b111100000000;
20'b01100101110110001111: color_data = 12'b111100000000;
20'b01100101110110010000: color_data = 12'b111100000000;
20'b01100101110110010001: color_data = 12'b111100000000;
20'b01100101110110010010: color_data = 12'b111100000000;
20'b01100101110110010011: color_data = 12'b111100000000;
20'b01100101110110010100: color_data = 12'b111100000000;
20'b01100101110110010101: color_data = 12'b111100000000;
20'b01100101110110010110: color_data = 12'b111100000000;
20'b01100101110110010111: color_data = 12'b111100000000;
20'b01100101110110011000: color_data = 12'b111100000000;
20'b01100101110110011001: color_data = 12'b111100000000;
20'b01100101110110011010: color_data = 12'b111100000000;
20'b01100101110110011011: color_data = 12'b111100000000;
20'b01100101110110011100: color_data = 12'b111100000000;
20'b01100101110110011101: color_data = 12'b111100000000;
20'b01100101110110011110: color_data = 12'b111100000000;
20'b01100110000011111010: color_data = 12'b000001101111;
20'b01100110000011111011: color_data = 12'b000001101111;
20'b01100110000011111100: color_data = 12'b000001101111;
20'b01100110000011111101: color_data = 12'b000001101111;
20'b01100110000011111110: color_data = 12'b000001101111;
20'b01100110000011111111: color_data = 12'b000001101111;
20'b01100110000100000000: color_data = 12'b000001101111;
20'b01100110000100000001: color_data = 12'b000001101111;
20'b01100110000100000010: color_data = 12'b000001101111;
20'b01100110000100000011: color_data = 12'b000001101111;
20'b01100110000100000100: color_data = 12'b000001101111;
20'b01100110000100000101: color_data = 12'b000001101111;
20'b01100110000100000110: color_data = 12'b000001101111;
20'b01100110000100000111: color_data = 12'b000001101111;
20'b01100110000100001000: color_data = 12'b000001101111;
20'b01100110000100001001: color_data = 12'b000001101111;
20'b01100110000100001010: color_data = 12'b000001101111;
20'b01100110000100001011: color_data = 12'b000001101111;
20'b01100110000100001111: color_data = 12'b000001101111;
20'b01100110000100010000: color_data = 12'b000001101111;
20'b01100110000100010001: color_data = 12'b000001101111;
20'b01100110000100010010: color_data = 12'b000001101111;
20'b01100110000100010011: color_data = 12'b000001101111;
20'b01100110000100010100: color_data = 12'b000001101111;
20'b01100110000100010101: color_data = 12'b000001101111;
20'b01100110000100010110: color_data = 12'b000001101111;
20'b01100110000100010111: color_data = 12'b000001101111;
20'b01100110000100011000: color_data = 12'b000001101111;
20'b01100110000100011001: color_data = 12'b000001101111;
20'b01100110000100011010: color_data = 12'b000001101111;
20'b01100110000100011011: color_data = 12'b000001101111;
20'b01100110000100011100: color_data = 12'b000001101111;
20'b01100110000100011101: color_data = 12'b000001101111;
20'b01100110000100011110: color_data = 12'b000001101111;
20'b01100110000100011111: color_data = 12'b000001101111;
20'b01100110000100100000: color_data = 12'b000001101111;
20'b01100110000100100100: color_data = 12'b000001101111;
20'b01100110000100100101: color_data = 12'b000001101111;
20'b01100110000100100110: color_data = 12'b000001101111;
20'b01100110000100100111: color_data = 12'b000001101111;
20'b01100110000100101000: color_data = 12'b000001101111;
20'b01100110000100101001: color_data = 12'b000001101111;
20'b01100110000100101010: color_data = 12'b000001101111;
20'b01100110000100101011: color_data = 12'b000001101111;
20'b01100110000100101100: color_data = 12'b000001101111;
20'b01100110000100101101: color_data = 12'b000001101111;
20'b01100110000100101110: color_data = 12'b000001101111;
20'b01100110000100101111: color_data = 12'b000001101111;
20'b01100110000100110000: color_data = 12'b000001101111;
20'b01100110000100110001: color_data = 12'b000001101111;
20'b01100110000100110010: color_data = 12'b000001101111;
20'b01100110000100110011: color_data = 12'b000001101111;
20'b01100110000100110100: color_data = 12'b000001101111;
20'b01100110000100110101: color_data = 12'b000001101111;
20'b01100110000100111001: color_data = 12'b000011110000;
20'b01100110000100111010: color_data = 12'b000011110000;
20'b01100110000100111011: color_data = 12'b000011110000;
20'b01100110000100111100: color_data = 12'b000011110000;
20'b01100110000100111101: color_data = 12'b000011110000;
20'b01100110000100111110: color_data = 12'b000011110000;
20'b01100110000100111111: color_data = 12'b000011110000;
20'b01100110000101000000: color_data = 12'b000011110000;
20'b01100110000101000001: color_data = 12'b000011110000;
20'b01100110000101000010: color_data = 12'b000011110000;
20'b01100110000101000011: color_data = 12'b000011110000;
20'b01100110000101000100: color_data = 12'b000011110000;
20'b01100110000101000101: color_data = 12'b000011110000;
20'b01100110000101000110: color_data = 12'b000011110000;
20'b01100110000101000111: color_data = 12'b000011110000;
20'b01100110000101001000: color_data = 12'b000011110000;
20'b01100110000101001001: color_data = 12'b000011110000;
20'b01100110000101001010: color_data = 12'b000011110000;
20'b01100110000101001110: color_data = 12'b000011110000;
20'b01100110000101001111: color_data = 12'b000011110000;
20'b01100110000101010000: color_data = 12'b000011110000;
20'b01100110000101010001: color_data = 12'b000011110000;
20'b01100110000101010010: color_data = 12'b000011110000;
20'b01100110000101010011: color_data = 12'b000011110000;
20'b01100110000101010100: color_data = 12'b000011110000;
20'b01100110000101010101: color_data = 12'b000011110000;
20'b01100110000101010110: color_data = 12'b000011110000;
20'b01100110000101010111: color_data = 12'b000011110000;
20'b01100110000101011000: color_data = 12'b000011110000;
20'b01100110000101011001: color_data = 12'b000011110000;
20'b01100110000101011010: color_data = 12'b000011110000;
20'b01100110000101011011: color_data = 12'b000011110000;
20'b01100110000101011100: color_data = 12'b000011110000;
20'b01100110000101011101: color_data = 12'b000011110000;
20'b01100110000101011110: color_data = 12'b000011110000;
20'b01100110000101011111: color_data = 12'b000011110000;
20'b01100110000101100011: color_data = 12'b111100001111;
20'b01100110000101100100: color_data = 12'b111100001111;
20'b01100110000101100101: color_data = 12'b111100001111;
20'b01100110000101100110: color_data = 12'b111100001111;
20'b01100110000101100111: color_data = 12'b111100001111;
20'b01100110000101101000: color_data = 12'b111100001111;
20'b01100110000101101001: color_data = 12'b111100001111;
20'b01100110000101101010: color_data = 12'b111100001111;
20'b01100110000101101011: color_data = 12'b111100001111;
20'b01100110000101101100: color_data = 12'b111100001111;
20'b01100110000101101101: color_data = 12'b111100001111;
20'b01100110000101101110: color_data = 12'b111100001111;
20'b01100110000101101111: color_data = 12'b111100001111;
20'b01100110000101110000: color_data = 12'b111100001111;
20'b01100110000101110001: color_data = 12'b111100001111;
20'b01100110000101110010: color_data = 12'b111100001111;
20'b01100110000101110011: color_data = 12'b111100001111;
20'b01100110000101110100: color_data = 12'b111100001111;
20'b01100110000101111000: color_data = 12'b111100001111;
20'b01100110000101111001: color_data = 12'b111100001111;
20'b01100110000101111010: color_data = 12'b111100001111;
20'b01100110000101111011: color_data = 12'b111100001111;
20'b01100110000101111100: color_data = 12'b111100001111;
20'b01100110000101111101: color_data = 12'b111100001111;
20'b01100110000101111110: color_data = 12'b111100001111;
20'b01100110000101111111: color_data = 12'b111100001111;
20'b01100110000110000000: color_data = 12'b111100001111;
20'b01100110000110000001: color_data = 12'b111100001111;
20'b01100110000110000010: color_data = 12'b111100001111;
20'b01100110000110000011: color_data = 12'b111100001111;
20'b01100110000110000100: color_data = 12'b111100001111;
20'b01100110000110000101: color_data = 12'b111100001111;
20'b01100110000110000110: color_data = 12'b111100001111;
20'b01100110000110000111: color_data = 12'b111100001111;
20'b01100110000110001000: color_data = 12'b111100001111;
20'b01100110000110001001: color_data = 12'b111100001111;
20'b01100110000110001101: color_data = 12'b111100000000;
20'b01100110000110001110: color_data = 12'b111100000000;
20'b01100110000110001111: color_data = 12'b111100000000;
20'b01100110000110010000: color_data = 12'b111100000000;
20'b01100110000110010001: color_data = 12'b111100000000;
20'b01100110000110010010: color_data = 12'b111100000000;
20'b01100110000110010011: color_data = 12'b111100000000;
20'b01100110000110010100: color_data = 12'b111100000000;
20'b01100110000110010101: color_data = 12'b111100000000;
20'b01100110000110010110: color_data = 12'b111100000000;
20'b01100110000110010111: color_data = 12'b111100000000;
20'b01100110000110011000: color_data = 12'b111100000000;
20'b01100110000110011001: color_data = 12'b111100000000;
20'b01100110000110011010: color_data = 12'b111100000000;
20'b01100110000110011011: color_data = 12'b111100000000;
20'b01100110000110011100: color_data = 12'b111100000000;
20'b01100110000110011101: color_data = 12'b111100000000;
20'b01100110000110011110: color_data = 12'b111100000000;
20'b01100110010011111010: color_data = 12'b000001101111;
20'b01100110010011111011: color_data = 12'b000001101111;
20'b01100110010011111100: color_data = 12'b000001101111;
20'b01100110010011111101: color_data = 12'b000001101111;
20'b01100110010011111110: color_data = 12'b000001101111;
20'b01100110010011111111: color_data = 12'b000001101111;
20'b01100110010100000000: color_data = 12'b000001101111;
20'b01100110010100000001: color_data = 12'b000001101111;
20'b01100110010100000010: color_data = 12'b000001101111;
20'b01100110010100000011: color_data = 12'b000001101111;
20'b01100110010100000100: color_data = 12'b000001101111;
20'b01100110010100000101: color_data = 12'b000001101111;
20'b01100110010100000110: color_data = 12'b000001101111;
20'b01100110010100000111: color_data = 12'b000001101111;
20'b01100110010100001000: color_data = 12'b000001101111;
20'b01100110010100001001: color_data = 12'b000001101111;
20'b01100110010100001010: color_data = 12'b000001101111;
20'b01100110010100001011: color_data = 12'b000001101111;
20'b01100110010100001111: color_data = 12'b000001101111;
20'b01100110010100010000: color_data = 12'b000001101111;
20'b01100110010100010001: color_data = 12'b000001101111;
20'b01100110010100010010: color_data = 12'b000001101111;
20'b01100110010100010011: color_data = 12'b000001101111;
20'b01100110010100010100: color_data = 12'b000001101111;
20'b01100110010100010101: color_data = 12'b000001101111;
20'b01100110010100010110: color_data = 12'b000001101111;
20'b01100110010100010111: color_data = 12'b000001101111;
20'b01100110010100011000: color_data = 12'b000001101111;
20'b01100110010100011001: color_data = 12'b000001101111;
20'b01100110010100011010: color_data = 12'b000001101111;
20'b01100110010100011011: color_data = 12'b000001101111;
20'b01100110010100011100: color_data = 12'b000001101111;
20'b01100110010100011101: color_data = 12'b000001101111;
20'b01100110010100011110: color_data = 12'b000001101111;
20'b01100110010100011111: color_data = 12'b000001101111;
20'b01100110010100100000: color_data = 12'b000001101111;
20'b01100110010100100100: color_data = 12'b000001101111;
20'b01100110010100100101: color_data = 12'b000001101111;
20'b01100110010100100110: color_data = 12'b000001101111;
20'b01100110010100100111: color_data = 12'b000001101111;
20'b01100110010100101000: color_data = 12'b000001101111;
20'b01100110010100101001: color_data = 12'b000001101111;
20'b01100110010100101010: color_data = 12'b000001101111;
20'b01100110010100101011: color_data = 12'b000001101111;
20'b01100110010100101100: color_data = 12'b000001101111;
20'b01100110010100101101: color_data = 12'b000001101111;
20'b01100110010100101110: color_data = 12'b000001101111;
20'b01100110010100101111: color_data = 12'b000001101111;
20'b01100110010100110000: color_data = 12'b000001101111;
20'b01100110010100110001: color_data = 12'b000001101111;
20'b01100110010100110010: color_data = 12'b000001101111;
20'b01100110010100110011: color_data = 12'b000001101111;
20'b01100110010100110100: color_data = 12'b000001101111;
20'b01100110010100110101: color_data = 12'b000001101111;
20'b01100110010100111001: color_data = 12'b000011110000;
20'b01100110010100111010: color_data = 12'b000011110000;
20'b01100110010100111011: color_data = 12'b000011110000;
20'b01100110010100111100: color_data = 12'b000011110000;
20'b01100110010100111101: color_data = 12'b000011110000;
20'b01100110010100111110: color_data = 12'b000011110000;
20'b01100110010100111111: color_data = 12'b000011110000;
20'b01100110010101000000: color_data = 12'b000011110000;
20'b01100110010101000001: color_data = 12'b000011110000;
20'b01100110010101000010: color_data = 12'b000011110000;
20'b01100110010101000011: color_data = 12'b000011110000;
20'b01100110010101000100: color_data = 12'b000011110000;
20'b01100110010101000101: color_data = 12'b000011110000;
20'b01100110010101000110: color_data = 12'b000011110000;
20'b01100110010101000111: color_data = 12'b000011110000;
20'b01100110010101001000: color_data = 12'b000011110000;
20'b01100110010101001001: color_data = 12'b000011110000;
20'b01100110010101001010: color_data = 12'b000011110000;
20'b01100110010101001110: color_data = 12'b000011110000;
20'b01100110010101001111: color_data = 12'b000011110000;
20'b01100110010101010000: color_data = 12'b000011110000;
20'b01100110010101010001: color_data = 12'b000011110000;
20'b01100110010101010010: color_data = 12'b000011110000;
20'b01100110010101010011: color_data = 12'b000011110000;
20'b01100110010101010100: color_data = 12'b000011110000;
20'b01100110010101010101: color_data = 12'b000011110000;
20'b01100110010101010110: color_data = 12'b000011110000;
20'b01100110010101010111: color_data = 12'b000011110000;
20'b01100110010101011000: color_data = 12'b000011110000;
20'b01100110010101011001: color_data = 12'b000011110000;
20'b01100110010101011010: color_data = 12'b000011110000;
20'b01100110010101011011: color_data = 12'b000011110000;
20'b01100110010101011100: color_data = 12'b000011110000;
20'b01100110010101011101: color_data = 12'b000011110000;
20'b01100110010101011110: color_data = 12'b000011110000;
20'b01100110010101011111: color_data = 12'b000011110000;
20'b01100110010101100011: color_data = 12'b111100001111;
20'b01100110010101100100: color_data = 12'b111100001111;
20'b01100110010101100101: color_data = 12'b111100001111;
20'b01100110010101100110: color_data = 12'b111100001111;
20'b01100110010101100111: color_data = 12'b111100001111;
20'b01100110010101101000: color_data = 12'b111100001111;
20'b01100110010101101001: color_data = 12'b111100001111;
20'b01100110010101101010: color_data = 12'b111100001111;
20'b01100110010101101011: color_data = 12'b111100001111;
20'b01100110010101101100: color_data = 12'b111100001111;
20'b01100110010101101101: color_data = 12'b111100001111;
20'b01100110010101101110: color_data = 12'b111100001111;
20'b01100110010101101111: color_data = 12'b111100001111;
20'b01100110010101110000: color_data = 12'b111100001111;
20'b01100110010101110001: color_data = 12'b111100001111;
20'b01100110010101110010: color_data = 12'b111100001111;
20'b01100110010101110011: color_data = 12'b111100001111;
20'b01100110010101110100: color_data = 12'b111100001111;
20'b01100110010101111000: color_data = 12'b111100001111;
20'b01100110010101111001: color_data = 12'b111100001111;
20'b01100110010101111010: color_data = 12'b111100001111;
20'b01100110010101111011: color_data = 12'b111100001111;
20'b01100110010101111100: color_data = 12'b111100001111;
20'b01100110010101111101: color_data = 12'b111100001111;
20'b01100110010101111110: color_data = 12'b111100001111;
20'b01100110010101111111: color_data = 12'b111100001111;
20'b01100110010110000000: color_data = 12'b111100001111;
20'b01100110010110000001: color_data = 12'b111100001111;
20'b01100110010110000010: color_data = 12'b111100001111;
20'b01100110010110000011: color_data = 12'b111100001111;
20'b01100110010110000100: color_data = 12'b111100001111;
20'b01100110010110000101: color_data = 12'b111100001111;
20'b01100110010110000110: color_data = 12'b111100001111;
20'b01100110010110000111: color_data = 12'b111100001111;
20'b01100110010110001000: color_data = 12'b111100001111;
20'b01100110010110001001: color_data = 12'b111100001111;
20'b01100110010110001101: color_data = 12'b111100000000;
20'b01100110010110001110: color_data = 12'b111100000000;
20'b01100110010110001111: color_data = 12'b111100000000;
20'b01100110010110010000: color_data = 12'b111100000000;
20'b01100110010110010001: color_data = 12'b111100000000;
20'b01100110010110010010: color_data = 12'b111100000000;
20'b01100110010110010011: color_data = 12'b111100000000;
20'b01100110010110010100: color_data = 12'b111100000000;
20'b01100110010110010101: color_data = 12'b111100000000;
20'b01100110010110010110: color_data = 12'b111100000000;
20'b01100110010110010111: color_data = 12'b111100000000;
20'b01100110010110011000: color_data = 12'b111100000000;
20'b01100110010110011001: color_data = 12'b111100000000;
20'b01100110010110011010: color_data = 12'b111100000000;
20'b01100110010110011011: color_data = 12'b111100000000;
20'b01100110010110011100: color_data = 12'b111100000000;
20'b01100110010110011101: color_data = 12'b111100000000;
20'b01100110010110011110: color_data = 12'b111100000000;
20'b01100110100011111010: color_data = 12'b000001101111;
20'b01100110100011111011: color_data = 12'b000001101111;
20'b01100110100011111100: color_data = 12'b000001101111;
20'b01100110100011111101: color_data = 12'b000001101111;
20'b01100110100011111110: color_data = 12'b000001101111;
20'b01100110100011111111: color_data = 12'b000001101111;
20'b01100110100100000000: color_data = 12'b000001101111;
20'b01100110100100000001: color_data = 12'b000001101111;
20'b01100110100100000010: color_data = 12'b000001101111;
20'b01100110100100000011: color_data = 12'b000001101111;
20'b01100110100100000100: color_data = 12'b000001101111;
20'b01100110100100000101: color_data = 12'b000001101111;
20'b01100110100100000110: color_data = 12'b000001101111;
20'b01100110100100000111: color_data = 12'b000001101111;
20'b01100110100100001000: color_data = 12'b000001101111;
20'b01100110100100001001: color_data = 12'b000001101111;
20'b01100110100100001010: color_data = 12'b000001101111;
20'b01100110100100001011: color_data = 12'b000001101111;
20'b01100110100100001111: color_data = 12'b000001101111;
20'b01100110100100010000: color_data = 12'b000001101111;
20'b01100110100100010001: color_data = 12'b000001101111;
20'b01100110100100010010: color_data = 12'b000001101111;
20'b01100110100100010011: color_data = 12'b000001101111;
20'b01100110100100010100: color_data = 12'b000001101111;
20'b01100110100100010101: color_data = 12'b000001101111;
20'b01100110100100010110: color_data = 12'b000001101111;
20'b01100110100100010111: color_data = 12'b000001101111;
20'b01100110100100011000: color_data = 12'b000001101111;
20'b01100110100100011001: color_data = 12'b000001101111;
20'b01100110100100011010: color_data = 12'b000001101111;
20'b01100110100100011011: color_data = 12'b000001101111;
20'b01100110100100011100: color_data = 12'b000001101111;
20'b01100110100100011101: color_data = 12'b000001101111;
20'b01100110100100011110: color_data = 12'b000001101111;
20'b01100110100100011111: color_data = 12'b000001101111;
20'b01100110100100100000: color_data = 12'b000001101111;
20'b01100110100100100100: color_data = 12'b000001101111;
20'b01100110100100100101: color_data = 12'b000001101111;
20'b01100110100100100110: color_data = 12'b000001101111;
20'b01100110100100100111: color_data = 12'b000001101111;
20'b01100110100100101000: color_data = 12'b000001101111;
20'b01100110100100101001: color_data = 12'b000001101111;
20'b01100110100100101010: color_data = 12'b000001101111;
20'b01100110100100101011: color_data = 12'b000001101111;
20'b01100110100100101100: color_data = 12'b000001101111;
20'b01100110100100101101: color_data = 12'b000001101111;
20'b01100110100100101110: color_data = 12'b000001101111;
20'b01100110100100101111: color_data = 12'b000001101111;
20'b01100110100100110000: color_data = 12'b000001101111;
20'b01100110100100110001: color_data = 12'b000001101111;
20'b01100110100100110010: color_data = 12'b000001101111;
20'b01100110100100110011: color_data = 12'b000001101111;
20'b01100110100100110100: color_data = 12'b000001101111;
20'b01100110100100110101: color_data = 12'b000001101111;
20'b01100110100100111001: color_data = 12'b000011110000;
20'b01100110100100111010: color_data = 12'b000011110000;
20'b01100110100100111011: color_data = 12'b000011110000;
20'b01100110100100111100: color_data = 12'b000011110000;
20'b01100110100100111101: color_data = 12'b000011110000;
20'b01100110100100111110: color_data = 12'b000011110000;
20'b01100110100100111111: color_data = 12'b000011110000;
20'b01100110100101000000: color_data = 12'b000011110000;
20'b01100110100101000001: color_data = 12'b000011110000;
20'b01100110100101000010: color_data = 12'b000011110000;
20'b01100110100101000011: color_data = 12'b000011110000;
20'b01100110100101000100: color_data = 12'b000011110000;
20'b01100110100101000101: color_data = 12'b000011110000;
20'b01100110100101000110: color_data = 12'b000011110000;
20'b01100110100101000111: color_data = 12'b000011110000;
20'b01100110100101001000: color_data = 12'b000011110000;
20'b01100110100101001001: color_data = 12'b000011110000;
20'b01100110100101001010: color_data = 12'b000011110000;
20'b01100110100101001110: color_data = 12'b000011110000;
20'b01100110100101001111: color_data = 12'b000011110000;
20'b01100110100101010000: color_data = 12'b000011110000;
20'b01100110100101010001: color_data = 12'b000011110000;
20'b01100110100101010010: color_data = 12'b000011110000;
20'b01100110100101010011: color_data = 12'b000011110000;
20'b01100110100101010100: color_data = 12'b000011110000;
20'b01100110100101010101: color_data = 12'b000011110000;
20'b01100110100101010110: color_data = 12'b000011110000;
20'b01100110100101010111: color_data = 12'b000011110000;
20'b01100110100101011000: color_data = 12'b000011110000;
20'b01100110100101011001: color_data = 12'b000011110000;
20'b01100110100101011010: color_data = 12'b000011110000;
20'b01100110100101011011: color_data = 12'b000011110000;
20'b01100110100101011100: color_data = 12'b000011110000;
20'b01100110100101011101: color_data = 12'b000011110000;
20'b01100110100101011110: color_data = 12'b000011110000;
20'b01100110100101011111: color_data = 12'b000011110000;
20'b01100110100101100011: color_data = 12'b111100001111;
20'b01100110100101100100: color_data = 12'b111100001111;
20'b01100110100101100101: color_data = 12'b111100001111;
20'b01100110100101100110: color_data = 12'b111100001111;
20'b01100110100101100111: color_data = 12'b111100001111;
20'b01100110100101101000: color_data = 12'b111100001111;
20'b01100110100101101001: color_data = 12'b111100001111;
20'b01100110100101101010: color_data = 12'b111100001111;
20'b01100110100101101011: color_data = 12'b111100001111;
20'b01100110100101101100: color_data = 12'b111100001111;
20'b01100110100101101101: color_data = 12'b111100001111;
20'b01100110100101101110: color_data = 12'b111100001111;
20'b01100110100101101111: color_data = 12'b111100001111;
20'b01100110100101110000: color_data = 12'b111100001111;
20'b01100110100101110001: color_data = 12'b111100001111;
20'b01100110100101110010: color_data = 12'b111100001111;
20'b01100110100101110011: color_data = 12'b111100001111;
20'b01100110100101110100: color_data = 12'b111100001111;
20'b01100110100101111000: color_data = 12'b111100001111;
20'b01100110100101111001: color_data = 12'b111100001111;
20'b01100110100101111010: color_data = 12'b111100001111;
20'b01100110100101111011: color_data = 12'b111100001111;
20'b01100110100101111100: color_data = 12'b111100001111;
20'b01100110100101111101: color_data = 12'b111100001111;
20'b01100110100101111110: color_data = 12'b111100001111;
20'b01100110100101111111: color_data = 12'b111100001111;
20'b01100110100110000000: color_data = 12'b111100001111;
20'b01100110100110000001: color_data = 12'b111100001111;
20'b01100110100110000010: color_data = 12'b111100001111;
20'b01100110100110000011: color_data = 12'b111100001111;
20'b01100110100110000100: color_data = 12'b111100001111;
20'b01100110100110000101: color_data = 12'b111100001111;
20'b01100110100110000110: color_data = 12'b111100001111;
20'b01100110100110000111: color_data = 12'b111100001111;
20'b01100110100110001000: color_data = 12'b111100001111;
20'b01100110100110001001: color_data = 12'b111100001111;
20'b01100110100110001101: color_data = 12'b111100000000;
20'b01100110100110001110: color_data = 12'b111100000000;
20'b01100110100110001111: color_data = 12'b111100000000;
20'b01100110100110010000: color_data = 12'b111100000000;
20'b01100110100110010001: color_data = 12'b111100000000;
20'b01100110100110010010: color_data = 12'b111100000000;
20'b01100110100110010011: color_data = 12'b111100000000;
20'b01100110100110010100: color_data = 12'b111100000000;
20'b01100110100110010101: color_data = 12'b111100000000;
20'b01100110100110010110: color_data = 12'b111100000000;
20'b01100110100110010111: color_data = 12'b111100000000;
20'b01100110100110011000: color_data = 12'b111100000000;
20'b01100110100110011001: color_data = 12'b111100000000;
20'b01100110100110011010: color_data = 12'b111100000000;
20'b01100110100110011011: color_data = 12'b111100000000;
20'b01100110100110011100: color_data = 12'b111100000000;
20'b01100110100110011101: color_data = 12'b111100000000;
20'b01100110100110011110: color_data = 12'b111100000000;
20'b01100110110011111010: color_data = 12'b000001101111;
20'b01100110110011111011: color_data = 12'b000001101111;
20'b01100110110011111100: color_data = 12'b000001101111;
20'b01100110110011111101: color_data = 12'b000001101111;
20'b01100110110011111110: color_data = 12'b000001101111;
20'b01100110110011111111: color_data = 12'b000001101111;
20'b01100110110100000000: color_data = 12'b000001101111;
20'b01100110110100000001: color_data = 12'b000001101111;
20'b01100110110100000010: color_data = 12'b000001101111;
20'b01100110110100000011: color_data = 12'b000001101111;
20'b01100110110100000100: color_data = 12'b000001101111;
20'b01100110110100000101: color_data = 12'b000001101111;
20'b01100110110100000110: color_data = 12'b000001101111;
20'b01100110110100000111: color_data = 12'b000001101111;
20'b01100110110100001000: color_data = 12'b000001101111;
20'b01100110110100001001: color_data = 12'b000001101111;
20'b01100110110100001010: color_data = 12'b000001101111;
20'b01100110110100001011: color_data = 12'b000001101111;
20'b01100110110100001111: color_data = 12'b000001101111;
20'b01100110110100010000: color_data = 12'b000001101111;
20'b01100110110100010001: color_data = 12'b000001101111;
20'b01100110110100010010: color_data = 12'b000001101111;
20'b01100110110100010011: color_data = 12'b000001101111;
20'b01100110110100010100: color_data = 12'b000001101111;
20'b01100110110100010101: color_data = 12'b000001101111;
20'b01100110110100010110: color_data = 12'b000001101111;
20'b01100110110100010111: color_data = 12'b000001101111;
20'b01100110110100011000: color_data = 12'b000001101111;
20'b01100110110100011001: color_data = 12'b000001101111;
20'b01100110110100011010: color_data = 12'b000001101111;
20'b01100110110100011011: color_data = 12'b000001101111;
20'b01100110110100011100: color_data = 12'b000001101111;
20'b01100110110100011101: color_data = 12'b000001101111;
20'b01100110110100011110: color_data = 12'b000001101111;
20'b01100110110100011111: color_data = 12'b000001101111;
20'b01100110110100100000: color_data = 12'b000001101111;
20'b01100110110100100100: color_data = 12'b000001101111;
20'b01100110110100100101: color_data = 12'b000001101111;
20'b01100110110100100110: color_data = 12'b000001101111;
20'b01100110110100100111: color_data = 12'b000001101111;
20'b01100110110100101000: color_data = 12'b000001101111;
20'b01100110110100101001: color_data = 12'b000001101111;
20'b01100110110100101010: color_data = 12'b000001101111;
20'b01100110110100101011: color_data = 12'b000001101111;
20'b01100110110100101100: color_data = 12'b000001101111;
20'b01100110110100101101: color_data = 12'b000001101111;
20'b01100110110100101110: color_data = 12'b000001101111;
20'b01100110110100101111: color_data = 12'b000001101111;
20'b01100110110100110000: color_data = 12'b000001101111;
20'b01100110110100110001: color_data = 12'b000001101111;
20'b01100110110100110010: color_data = 12'b000001101111;
20'b01100110110100110011: color_data = 12'b000001101111;
20'b01100110110100110100: color_data = 12'b000001101111;
20'b01100110110100110101: color_data = 12'b000001101111;
20'b01100110110100111001: color_data = 12'b000011110000;
20'b01100110110100111010: color_data = 12'b000011110000;
20'b01100110110100111011: color_data = 12'b000011110000;
20'b01100110110100111100: color_data = 12'b000011110000;
20'b01100110110100111101: color_data = 12'b000011110000;
20'b01100110110100111110: color_data = 12'b000011110000;
20'b01100110110100111111: color_data = 12'b000011110000;
20'b01100110110101000000: color_data = 12'b000011110000;
20'b01100110110101000001: color_data = 12'b000011110000;
20'b01100110110101000010: color_data = 12'b000011110000;
20'b01100110110101000011: color_data = 12'b000011110000;
20'b01100110110101000100: color_data = 12'b000011110000;
20'b01100110110101000101: color_data = 12'b000011110000;
20'b01100110110101000110: color_data = 12'b000011110000;
20'b01100110110101000111: color_data = 12'b000011110000;
20'b01100110110101001000: color_data = 12'b000011110000;
20'b01100110110101001001: color_data = 12'b000011110000;
20'b01100110110101001010: color_data = 12'b000011110000;
20'b01100110110101001110: color_data = 12'b000011110000;
20'b01100110110101001111: color_data = 12'b000011110000;
20'b01100110110101010000: color_data = 12'b000011110000;
20'b01100110110101010001: color_data = 12'b000011110000;
20'b01100110110101010010: color_data = 12'b000011110000;
20'b01100110110101010011: color_data = 12'b000011110000;
20'b01100110110101010100: color_data = 12'b000011110000;
20'b01100110110101010101: color_data = 12'b000011110000;
20'b01100110110101010110: color_data = 12'b000011110000;
20'b01100110110101010111: color_data = 12'b000011110000;
20'b01100110110101011000: color_data = 12'b000011110000;
20'b01100110110101011001: color_data = 12'b000011110000;
20'b01100110110101011010: color_data = 12'b000011110000;
20'b01100110110101011011: color_data = 12'b000011110000;
20'b01100110110101011100: color_data = 12'b000011110000;
20'b01100110110101011101: color_data = 12'b000011110000;
20'b01100110110101011110: color_data = 12'b000011110000;
20'b01100110110101011111: color_data = 12'b000011110000;
20'b01100110110101100011: color_data = 12'b111100001111;
20'b01100110110101100100: color_data = 12'b111100001111;
20'b01100110110101100101: color_data = 12'b111100001111;
20'b01100110110101100110: color_data = 12'b111100001111;
20'b01100110110101100111: color_data = 12'b111100001111;
20'b01100110110101101000: color_data = 12'b111100001111;
20'b01100110110101101001: color_data = 12'b111100001111;
20'b01100110110101101010: color_data = 12'b111100001111;
20'b01100110110101101011: color_data = 12'b111100001111;
20'b01100110110101101100: color_data = 12'b111100001111;
20'b01100110110101101101: color_data = 12'b111100001111;
20'b01100110110101101110: color_data = 12'b111100001111;
20'b01100110110101101111: color_data = 12'b111100001111;
20'b01100110110101110000: color_data = 12'b111100001111;
20'b01100110110101110001: color_data = 12'b111100001111;
20'b01100110110101110010: color_data = 12'b111100001111;
20'b01100110110101110011: color_data = 12'b111100001111;
20'b01100110110101110100: color_data = 12'b111100001111;
20'b01100110110101111000: color_data = 12'b111100001111;
20'b01100110110101111001: color_data = 12'b111100001111;
20'b01100110110101111010: color_data = 12'b111100001111;
20'b01100110110101111011: color_data = 12'b111100001111;
20'b01100110110101111100: color_data = 12'b111100001111;
20'b01100110110101111101: color_data = 12'b111100001111;
20'b01100110110101111110: color_data = 12'b111100001111;
20'b01100110110101111111: color_data = 12'b111100001111;
20'b01100110110110000000: color_data = 12'b111100001111;
20'b01100110110110000001: color_data = 12'b111100001111;
20'b01100110110110000010: color_data = 12'b111100001111;
20'b01100110110110000011: color_data = 12'b111100001111;
20'b01100110110110000100: color_data = 12'b111100001111;
20'b01100110110110000101: color_data = 12'b111100001111;
20'b01100110110110000110: color_data = 12'b111100001111;
20'b01100110110110000111: color_data = 12'b111100001111;
20'b01100110110110001000: color_data = 12'b111100001111;
20'b01100110110110001001: color_data = 12'b111100001111;
20'b01100110110110001101: color_data = 12'b111100000000;
20'b01100110110110001110: color_data = 12'b111100000000;
20'b01100110110110001111: color_data = 12'b111100000000;
20'b01100110110110010000: color_data = 12'b111100000000;
20'b01100110110110010001: color_data = 12'b111100000000;
20'b01100110110110010010: color_data = 12'b111100000000;
20'b01100110110110010011: color_data = 12'b111100000000;
20'b01100110110110010100: color_data = 12'b111100000000;
20'b01100110110110010101: color_data = 12'b111100000000;
20'b01100110110110010110: color_data = 12'b111100000000;
20'b01100110110110010111: color_data = 12'b111100000000;
20'b01100110110110011000: color_data = 12'b111100000000;
20'b01100110110110011001: color_data = 12'b111100000000;
20'b01100110110110011010: color_data = 12'b111100000000;
20'b01100110110110011011: color_data = 12'b111100000000;
20'b01100110110110011100: color_data = 12'b111100000000;
20'b01100110110110011101: color_data = 12'b111100000000;
20'b01100110110110011110: color_data = 12'b111100000000;
20'b01100111000011111010: color_data = 12'b000001101111;
20'b01100111000011111011: color_data = 12'b000001101111;
20'b01100111000011111100: color_data = 12'b000001101111;
20'b01100111000011111101: color_data = 12'b000001101111;
20'b01100111000011111110: color_data = 12'b000001101111;
20'b01100111000011111111: color_data = 12'b000001101111;
20'b01100111000100000000: color_data = 12'b000001101111;
20'b01100111000100000001: color_data = 12'b000001101111;
20'b01100111000100000010: color_data = 12'b000001101111;
20'b01100111000100000011: color_data = 12'b000001101111;
20'b01100111000100000100: color_data = 12'b000001101111;
20'b01100111000100000101: color_data = 12'b000001101111;
20'b01100111000100000110: color_data = 12'b000001101111;
20'b01100111000100000111: color_data = 12'b000001101111;
20'b01100111000100001000: color_data = 12'b000001101111;
20'b01100111000100001001: color_data = 12'b000001101111;
20'b01100111000100001010: color_data = 12'b000001101111;
20'b01100111000100001011: color_data = 12'b000001101111;
20'b01100111000100001111: color_data = 12'b000001101111;
20'b01100111000100010000: color_data = 12'b000001101111;
20'b01100111000100010001: color_data = 12'b000001101111;
20'b01100111000100010010: color_data = 12'b000001101111;
20'b01100111000100010011: color_data = 12'b000001101111;
20'b01100111000100010100: color_data = 12'b000001101111;
20'b01100111000100010101: color_data = 12'b000001101111;
20'b01100111000100010110: color_data = 12'b000001101111;
20'b01100111000100010111: color_data = 12'b000001101111;
20'b01100111000100011000: color_data = 12'b000001101111;
20'b01100111000100011001: color_data = 12'b000001101111;
20'b01100111000100011010: color_data = 12'b000001101111;
20'b01100111000100011011: color_data = 12'b000001101111;
20'b01100111000100011100: color_data = 12'b000001101111;
20'b01100111000100011101: color_data = 12'b000001101111;
20'b01100111000100011110: color_data = 12'b000001101111;
20'b01100111000100011111: color_data = 12'b000001101111;
20'b01100111000100100000: color_data = 12'b000001101111;
20'b01100111000100100100: color_data = 12'b000001101111;
20'b01100111000100100101: color_data = 12'b000001101111;
20'b01100111000100100110: color_data = 12'b000001101111;
20'b01100111000100100111: color_data = 12'b000001101111;
20'b01100111000100101000: color_data = 12'b000001101111;
20'b01100111000100101001: color_data = 12'b000001101111;
20'b01100111000100101010: color_data = 12'b000001101111;
20'b01100111000100101011: color_data = 12'b000001101111;
20'b01100111000100101100: color_data = 12'b000001101111;
20'b01100111000100101101: color_data = 12'b000001101111;
20'b01100111000100101110: color_data = 12'b000001101111;
20'b01100111000100101111: color_data = 12'b000001101111;
20'b01100111000100110000: color_data = 12'b000001101111;
20'b01100111000100110001: color_data = 12'b000001101111;
20'b01100111000100110010: color_data = 12'b000001101111;
20'b01100111000100110011: color_data = 12'b000001101111;
20'b01100111000100110100: color_data = 12'b000001101111;
20'b01100111000100110101: color_data = 12'b000001101111;
20'b01100111000100111001: color_data = 12'b000011110000;
20'b01100111000100111010: color_data = 12'b000011110000;
20'b01100111000100111011: color_data = 12'b000011110000;
20'b01100111000100111100: color_data = 12'b000011110000;
20'b01100111000100111101: color_data = 12'b000011110000;
20'b01100111000100111110: color_data = 12'b000011110000;
20'b01100111000100111111: color_data = 12'b000011110000;
20'b01100111000101000000: color_data = 12'b000011110000;
20'b01100111000101000001: color_data = 12'b000011110000;
20'b01100111000101000010: color_data = 12'b000011110000;
20'b01100111000101000011: color_data = 12'b000011110000;
20'b01100111000101000100: color_data = 12'b000011110000;
20'b01100111000101000101: color_data = 12'b000011110000;
20'b01100111000101000110: color_data = 12'b000011110000;
20'b01100111000101000111: color_data = 12'b000011110000;
20'b01100111000101001000: color_data = 12'b000011110000;
20'b01100111000101001001: color_data = 12'b000011110000;
20'b01100111000101001010: color_data = 12'b000011110000;
20'b01100111000101001110: color_data = 12'b000011110000;
20'b01100111000101001111: color_data = 12'b000011110000;
20'b01100111000101010000: color_data = 12'b000011110000;
20'b01100111000101010001: color_data = 12'b000011110000;
20'b01100111000101010010: color_data = 12'b000011110000;
20'b01100111000101010011: color_data = 12'b000011110000;
20'b01100111000101010100: color_data = 12'b000011110000;
20'b01100111000101010101: color_data = 12'b000011110000;
20'b01100111000101010110: color_data = 12'b000011110000;
20'b01100111000101010111: color_data = 12'b000011110000;
20'b01100111000101011000: color_data = 12'b000011110000;
20'b01100111000101011001: color_data = 12'b000011110000;
20'b01100111000101011010: color_data = 12'b000011110000;
20'b01100111000101011011: color_data = 12'b000011110000;
20'b01100111000101011100: color_data = 12'b000011110000;
20'b01100111000101011101: color_data = 12'b000011110000;
20'b01100111000101011110: color_data = 12'b000011110000;
20'b01100111000101011111: color_data = 12'b000011110000;
20'b01100111000101100011: color_data = 12'b111100001111;
20'b01100111000101100100: color_data = 12'b111100001111;
20'b01100111000101100101: color_data = 12'b111100001111;
20'b01100111000101100110: color_data = 12'b111100001111;
20'b01100111000101100111: color_data = 12'b111100001111;
20'b01100111000101101000: color_data = 12'b111100001111;
20'b01100111000101101001: color_data = 12'b111100001111;
20'b01100111000101101010: color_data = 12'b111100001111;
20'b01100111000101101011: color_data = 12'b111100001111;
20'b01100111000101101100: color_data = 12'b111100001111;
20'b01100111000101101101: color_data = 12'b111100001111;
20'b01100111000101101110: color_data = 12'b111100001111;
20'b01100111000101101111: color_data = 12'b111100001111;
20'b01100111000101110000: color_data = 12'b111100001111;
20'b01100111000101110001: color_data = 12'b111100001111;
20'b01100111000101110010: color_data = 12'b111100001111;
20'b01100111000101110011: color_data = 12'b111100001111;
20'b01100111000101110100: color_data = 12'b111100001111;
20'b01100111000101111000: color_data = 12'b111100001111;
20'b01100111000101111001: color_data = 12'b111100001111;
20'b01100111000101111010: color_data = 12'b111100001111;
20'b01100111000101111011: color_data = 12'b111100001111;
20'b01100111000101111100: color_data = 12'b111100001111;
20'b01100111000101111101: color_data = 12'b111100001111;
20'b01100111000101111110: color_data = 12'b111100001111;
20'b01100111000101111111: color_data = 12'b111100001111;
20'b01100111000110000000: color_data = 12'b111100001111;
20'b01100111000110000001: color_data = 12'b111100001111;
20'b01100111000110000010: color_data = 12'b111100001111;
20'b01100111000110000011: color_data = 12'b111100001111;
20'b01100111000110000100: color_data = 12'b111100001111;
20'b01100111000110000101: color_data = 12'b111100001111;
20'b01100111000110000110: color_data = 12'b111100001111;
20'b01100111000110000111: color_data = 12'b111100001111;
20'b01100111000110001000: color_data = 12'b111100001111;
20'b01100111000110001001: color_data = 12'b111100001111;
20'b01100111000110001101: color_data = 12'b111100000000;
20'b01100111000110001110: color_data = 12'b111100000000;
20'b01100111000110001111: color_data = 12'b111100000000;
20'b01100111000110010000: color_data = 12'b111100000000;
20'b01100111000110010001: color_data = 12'b111100000000;
20'b01100111000110010010: color_data = 12'b111100000000;
20'b01100111000110010011: color_data = 12'b111100000000;
20'b01100111000110010100: color_data = 12'b111100000000;
20'b01100111000110010101: color_data = 12'b111100000000;
20'b01100111000110010110: color_data = 12'b111100000000;
20'b01100111000110010111: color_data = 12'b111100000000;
20'b01100111000110011000: color_data = 12'b111100000000;
20'b01100111000110011001: color_data = 12'b111100000000;
20'b01100111000110011010: color_data = 12'b111100000000;
20'b01100111000110011011: color_data = 12'b111100000000;
20'b01100111000110011100: color_data = 12'b111100000000;
20'b01100111000110011101: color_data = 12'b111100000000;
20'b01100111000110011110: color_data = 12'b111100000000;
20'b01100111010011111010: color_data = 12'b000001101111;
20'b01100111010011111011: color_data = 12'b000001101111;
20'b01100111010011111100: color_data = 12'b000001101111;
20'b01100111010011111101: color_data = 12'b000001101111;
20'b01100111010011111110: color_data = 12'b000001101111;
20'b01100111010011111111: color_data = 12'b000001101111;
20'b01100111010100000000: color_data = 12'b000001101111;
20'b01100111010100000001: color_data = 12'b000001101111;
20'b01100111010100000010: color_data = 12'b000001101111;
20'b01100111010100000011: color_data = 12'b000001101111;
20'b01100111010100000100: color_data = 12'b000001101111;
20'b01100111010100000101: color_data = 12'b000001101111;
20'b01100111010100000110: color_data = 12'b000001101111;
20'b01100111010100000111: color_data = 12'b000001101111;
20'b01100111010100001000: color_data = 12'b000001101111;
20'b01100111010100001001: color_data = 12'b000001101111;
20'b01100111010100001010: color_data = 12'b000001101111;
20'b01100111010100001011: color_data = 12'b000001101111;
20'b01100111010100001111: color_data = 12'b000001101111;
20'b01100111010100010000: color_data = 12'b000001101111;
20'b01100111010100010001: color_data = 12'b000001101111;
20'b01100111010100010010: color_data = 12'b000001101111;
20'b01100111010100010011: color_data = 12'b000001101111;
20'b01100111010100010100: color_data = 12'b000001101111;
20'b01100111010100010101: color_data = 12'b000001101111;
20'b01100111010100010110: color_data = 12'b000001101111;
20'b01100111010100010111: color_data = 12'b000001101111;
20'b01100111010100011000: color_data = 12'b000001101111;
20'b01100111010100011001: color_data = 12'b000001101111;
20'b01100111010100011010: color_data = 12'b000001101111;
20'b01100111010100011011: color_data = 12'b000001101111;
20'b01100111010100011100: color_data = 12'b000001101111;
20'b01100111010100011101: color_data = 12'b000001101111;
20'b01100111010100011110: color_data = 12'b000001101111;
20'b01100111010100011111: color_data = 12'b000001101111;
20'b01100111010100100000: color_data = 12'b000001101111;
20'b01100111010100100100: color_data = 12'b000001101111;
20'b01100111010100100101: color_data = 12'b000001101111;
20'b01100111010100100110: color_data = 12'b000001101111;
20'b01100111010100100111: color_data = 12'b000001101111;
20'b01100111010100101000: color_data = 12'b000001101111;
20'b01100111010100101001: color_data = 12'b000001101111;
20'b01100111010100101010: color_data = 12'b000001101111;
20'b01100111010100101011: color_data = 12'b000001101111;
20'b01100111010100101100: color_data = 12'b000001101111;
20'b01100111010100101101: color_data = 12'b000001101111;
20'b01100111010100101110: color_data = 12'b000001101111;
20'b01100111010100101111: color_data = 12'b000001101111;
20'b01100111010100110000: color_data = 12'b000001101111;
20'b01100111010100110001: color_data = 12'b000001101111;
20'b01100111010100110010: color_data = 12'b000001101111;
20'b01100111010100110011: color_data = 12'b000001101111;
20'b01100111010100110100: color_data = 12'b000001101111;
20'b01100111010100110101: color_data = 12'b000001101111;
20'b01100111010100111001: color_data = 12'b000011110000;
20'b01100111010100111010: color_data = 12'b000011110000;
20'b01100111010100111011: color_data = 12'b000011110000;
20'b01100111010100111100: color_data = 12'b000011110000;
20'b01100111010100111101: color_data = 12'b000011110000;
20'b01100111010100111110: color_data = 12'b000011110000;
20'b01100111010100111111: color_data = 12'b000011110000;
20'b01100111010101000000: color_data = 12'b000011110000;
20'b01100111010101000001: color_data = 12'b000011110000;
20'b01100111010101000010: color_data = 12'b000011110000;
20'b01100111010101000011: color_data = 12'b000011110000;
20'b01100111010101000100: color_data = 12'b000011110000;
20'b01100111010101000101: color_data = 12'b000011110000;
20'b01100111010101000110: color_data = 12'b000011110000;
20'b01100111010101000111: color_data = 12'b000011110000;
20'b01100111010101001000: color_data = 12'b000011110000;
20'b01100111010101001001: color_data = 12'b000011110000;
20'b01100111010101001010: color_data = 12'b000011110000;
20'b01100111010101001110: color_data = 12'b000011110000;
20'b01100111010101001111: color_data = 12'b000011110000;
20'b01100111010101010000: color_data = 12'b000011110000;
20'b01100111010101010001: color_data = 12'b000011110000;
20'b01100111010101010010: color_data = 12'b000011110000;
20'b01100111010101010011: color_data = 12'b000011110000;
20'b01100111010101010100: color_data = 12'b000011110000;
20'b01100111010101010101: color_data = 12'b000011110000;
20'b01100111010101010110: color_data = 12'b000011110000;
20'b01100111010101010111: color_data = 12'b000011110000;
20'b01100111010101011000: color_data = 12'b000011110000;
20'b01100111010101011001: color_data = 12'b000011110000;
20'b01100111010101011010: color_data = 12'b000011110000;
20'b01100111010101011011: color_data = 12'b000011110000;
20'b01100111010101011100: color_data = 12'b000011110000;
20'b01100111010101011101: color_data = 12'b000011110000;
20'b01100111010101011110: color_data = 12'b000011110000;
20'b01100111010101011111: color_data = 12'b000011110000;
20'b01100111010101100011: color_data = 12'b111100001111;
20'b01100111010101100100: color_data = 12'b111100001111;
20'b01100111010101100101: color_data = 12'b111100001111;
20'b01100111010101100110: color_data = 12'b111100001111;
20'b01100111010101100111: color_data = 12'b111100001111;
20'b01100111010101101000: color_data = 12'b111100001111;
20'b01100111010101101001: color_data = 12'b111100001111;
20'b01100111010101101010: color_data = 12'b111100001111;
20'b01100111010101101011: color_data = 12'b111100001111;
20'b01100111010101101100: color_data = 12'b111100001111;
20'b01100111010101101101: color_data = 12'b111100001111;
20'b01100111010101101110: color_data = 12'b111100001111;
20'b01100111010101101111: color_data = 12'b111100001111;
20'b01100111010101110000: color_data = 12'b111100001111;
20'b01100111010101110001: color_data = 12'b111100001111;
20'b01100111010101110010: color_data = 12'b111100001111;
20'b01100111010101110011: color_data = 12'b111100001111;
20'b01100111010101110100: color_data = 12'b111100001111;
20'b01100111010101111000: color_data = 12'b111100001111;
20'b01100111010101111001: color_data = 12'b111100001111;
20'b01100111010101111010: color_data = 12'b111100001111;
20'b01100111010101111011: color_data = 12'b111100001111;
20'b01100111010101111100: color_data = 12'b111100001111;
20'b01100111010101111101: color_data = 12'b111100001111;
20'b01100111010101111110: color_data = 12'b111100001111;
20'b01100111010101111111: color_data = 12'b111100001111;
20'b01100111010110000000: color_data = 12'b111100001111;
20'b01100111010110000001: color_data = 12'b111100001111;
20'b01100111010110000010: color_data = 12'b111100001111;
20'b01100111010110000011: color_data = 12'b111100001111;
20'b01100111010110000100: color_data = 12'b111100001111;
20'b01100111010110000101: color_data = 12'b111100001111;
20'b01100111010110000110: color_data = 12'b111100001111;
20'b01100111010110000111: color_data = 12'b111100001111;
20'b01100111010110001000: color_data = 12'b111100001111;
20'b01100111010110001001: color_data = 12'b111100001111;
20'b01100111010110001101: color_data = 12'b111100000000;
20'b01100111010110001110: color_data = 12'b111100000000;
20'b01100111010110001111: color_data = 12'b111100000000;
20'b01100111010110010000: color_data = 12'b111100000000;
20'b01100111010110010001: color_data = 12'b111100000000;
20'b01100111010110010010: color_data = 12'b111100000000;
20'b01100111010110010011: color_data = 12'b111100000000;
20'b01100111010110010100: color_data = 12'b111100000000;
20'b01100111010110010101: color_data = 12'b111100000000;
20'b01100111010110010110: color_data = 12'b111100000000;
20'b01100111010110010111: color_data = 12'b111100000000;
20'b01100111010110011000: color_data = 12'b111100000000;
20'b01100111010110011001: color_data = 12'b111100000000;
20'b01100111010110011010: color_data = 12'b111100000000;
20'b01100111010110011011: color_data = 12'b111100000000;
20'b01100111010110011100: color_data = 12'b111100000000;
20'b01100111010110011101: color_data = 12'b111100000000;
20'b01100111010110011110: color_data = 12'b111100000000;
20'b01100111100011111010: color_data = 12'b000001101111;
20'b01100111100011111011: color_data = 12'b000001101111;
20'b01100111100011111100: color_data = 12'b000001101111;
20'b01100111100011111101: color_data = 12'b000001101111;
20'b01100111100011111110: color_data = 12'b000001101111;
20'b01100111100011111111: color_data = 12'b000001101111;
20'b01100111100100000000: color_data = 12'b000001101111;
20'b01100111100100000001: color_data = 12'b000001101111;
20'b01100111100100000010: color_data = 12'b000001101111;
20'b01100111100100000011: color_data = 12'b000001101111;
20'b01100111100100000100: color_data = 12'b000001101111;
20'b01100111100100000101: color_data = 12'b000001101111;
20'b01100111100100000110: color_data = 12'b000001101111;
20'b01100111100100000111: color_data = 12'b000001101111;
20'b01100111100100001000: color_data = 12'b000001101111;
20'b01100111100100001001: color_data = 12'b000001101111;
20'b01100111100100001010: color_data = 12'b000001101111;
20'b01100111100100001011: color_data = 12'b000001101111;
20'b01100111100100001111: color_data = 12'b000001101111;
20'b01100111100100010000: color_data = 12'b000001101111;
20'b01100111100100010001: color_data = 12'b000001101111;
20'b01100111100100010010: color_data = 12'b000001101111;
20'b01100111100100010011: color_data = 12'b000001101111;
20'b01100111100100010100: color_data = 12'b000001101111;
20'b01100111100100010101: color_data = 12'b000001101111;
20'b01100111100100010110: color_data = 12'b000001101111;
20'b01100111100100010111: color_data = 12'b000001101111;
20'b01100111100100011000: color_data = 12'b000001101111;
20'b01100111100100011001: color_data = 12'b000001101111;
20'b01100111100100011010: color_data = 12'b000001101111;
20'b01100111100100011011: color_data = 12'b000001101111;
20'b01100111100100011100: color_data = 12'b000001101111;
20'b01100111100100011101: color_data = 12'b000001101111;
20'b01100111100100011110: color_data = 12'b000001101111;
20'b01100111100100011111: color_data = 12'b000001101111;
20'b01100111100100100000: color_data = 12'b000001101111;
20'b01100111100100100100: color_data = 12'b000001101111;
20'b01100111100100100101: color_data = 12'b000001101111;
20'b01100111100100100110: color_data = 12'b000001101111;
20'b01100111100100100111: color_data = 12'b000001101111;
20'b01100111100100101000: color_data = 12'b000001101111;
20'b01100111100100101001: color_data = 12'b000001101111;
20'b01100111100100101010: color_data = 12'b000001101111;
20'b01100111100100101011: color_data = 12'b000001101111;
20'b01100111100100101100: color_data = 12'b000001101111;
20'b01100111100100101101: color_data = 12'b000001101111;
20'b01100111100100101110: color_data = 12'b000001101111;
20'b01100111100100101111: color_data = 12'b000001101111;
20'b01100111100100110000: color_data = 12'b000001101111;
20'b01100111100100110001: color_data = 12'b000001101111;
20'b01100111100100110010: color_data = 12'b000001101111;
20'b01100111100100110011: color_data = 12'b000001101111;
20'b01100111100100110100: color_data = 12'b000001101111;
20'b01100111100100110101: color_data = 12'b000001101111;
20'b01100111100100111001: color_data = 12'b000011110000;
20'b01100111100100111010: color_data = 12'b000011110000;
20'b01100111100100111011: color_data = 12'b000011110000;
20'b01100111100100111100: color_data = 12'b000011110000;
20'b01100111100100111101: color_data = 12'b000011110000;
20'b01100111100100111110: color_data = 12'b000011110000;
20'b01100111100100111111: color_data = 12'b000011110000;
20'b01100111100101000000: color_data = 12'b000011110000;
20'b01100111100101000001: color_data = 12'b000011110000;
20'b01100111100101000010: color_data = 12'b000011110000;
20'b01100111100101000011: color_data = 12'b000011110000;
20'b01100111100101000100: color_data = 12'b000011110000;
20'b01100111100101000101: color_data = 12'b000011110000;
20'b01100111100101000110: color_data = 12'b000011110000;
20'b01100111100101000111: color_data = 12'b000011110000;
20'b01100111100101001000: color_data = 12'b000011110000;
20'b01100111100101001001: color_data = 12'b000011110000;
20'b01100111100101001010: color_data = 12'b000011110000;
20'b01100111100101001110: color_data = 12'b000011110000;
20'b01100111100101001111: color_data = 12'b000011110000;
20'b01100111100101010000: color_data = 12'b000011110000;
20'b01100111100101010001: color_data = 12'b000011110000;
20'b01100111100101010010: color_data = 12'b000011110000;
20'b01100111100101010011: color_data = 12'b000011110000;
20'b01100111100101010100: color_data = 12'b000011110000;
20'b01100111100101010101: color_data = 12'b000011110000;
20'b01100111100101010110: color_data = 12'b000011110000;
20'b01100111100101010111: color_data = 12'b000011110000;
20'b01100111100101011000: color_data = 12'b000011110000;
20'b01100111100101011001: color_data = 12'b000011110000;
20'b01100111100101011010: color_data = 12'b000011110000;
20'b01100111100101011011: color_data = 12'b000011110000;
20'b01100111100101011100: color_data = 12'b000011110000;
20'b01100111100101011101: color_data = 12'b000011110000;
20'b01100111100101011110: color_data = 12'b000011110000;
20'b01100111100101011111: color_data = 12'b000011110000;
20'b01100111100101100011: color_data = 12'b111100001111;
20'b01100111100101100100: color_data = 12'b111100001111;
20'b01100111100101100101: color_data = 12'b111100001111;
20'b01100111100101100110: color_data = 12'b111100001111;
20'b01100111100101100111: color_data = 12'b111100001111;
20'b01100111100101101000: color_data = 12'b111100001111;
20'b01100111100101101001: color_data = 12'b111100001111;
20'b01100111100101101010: color_data = 12'b111100001111;
20'b01100111100101101011: color_data = 12'b111100001111;
20'b01100111100101101100: color_data = 12'b111100001111;
20'b01100111100101101101: color_data = 12'b111100001111;
20'b01100111100101101110: color_data = 12'b111100001111;
20'b01100111100101101111: color_data = 12'b111100001111;
20'b01100111100101110000: color_data = 12'b111100001111;
20'b01100111100101110001: color_data = 12'b111100001111;
20'b01100111100101110010: color_data = 12'b111100001111;
20'b01100111100101110011: color_data = 12'b111100001111;
20'b01100111100101110100: color_data = 12'b111100001111;
20'b01100111100101111000: color_data = 12'b111100001111;
20'b01100111100101111001: color_data = 12'b111100001111;
20'b01100111100101111010: color_data = 12'b111100001111;
20'b01100111100101111011: color_data = 12'b111100001111;
20'b01100111100101111100: color_data = 12'b111100001111;
20'b01100111100101111101: color_data = 12'b111100001111;
20'b01100111100101111110: color_data = 12'b111100001111;
20'b01100111100101111111: color_data = 12'b111100001111;
20'b01100111100110000000: color_data = 12'b111100001111;
20'b01100111100110000001: color_data = 12'b111100001111;
20'b01100111100110000010: color_data = 12'b111100001111;
20'b01100111100110000011: color_data = 12'b111100001111;
20'b01100111100110000100: color_data = 12'b111100001111;
20'b01100111100110000101: color_data = 12'b111100001111;
20'b01100111100110000110: color_data = 12'b111100001111;
20'b01100111100110000111: color_data = 12'b111100001111;
20'b01100111100110001000: color_data = 12'b111100001111;
20'b01100111100110001001: color_data = 12'b111100001111;
20'b01100111100110001101: color_data = 12'b111100000000;
20'b01100111100110001110: color_data = 12'b111100000000;
20'b01100111100110001111: color_data = 12'b111100000000;
20'b01100111100110010000: color_data = 12'b111100000000;
20'b01100111100110010001: color_data = 12'b111100000000;
20'b01100111100110010010: color_data = 12'b111100000000;
20'b01100111100110010011: color_data = 12'b111100000000;
20'b01100111100110010100: color_data = 12'b111100000000;
20'b01100111100110010101: color_data = 12'b111100000000;
20'b01100111100110010110: color_data = 12'b111100000000;
20'b01100111100110010111: color_data = 12'b111100000000;
20'b01100111100110011000: color_data = 12'b111100000000;
20'b01100111100110011001: color_data = 12'b111100000000;
20'b01100111100110011010: color_data = 12'b111100000000;
20'b01100111100110011011: color_data = 12'b111100000000;
20'b01100111100110011100: color_data = 12'b111100000000;
20'b01100111100110011101: color_data = 12'b111100000000;
20'b01100111100110011110: color_data = 12'b111100000000;
20'b01100111110011111010: color_data = 12'b000001101111;
20'b01100111110011111011: color_data = 12'b000001101111;
20'b01100111110011111100: color_data = 12'b000001101111;
20'b01100111110011111101: color_data = 12'b000001101111;
20'b01100111110011111110: color_data = 12'b000001101111;
20'b01100111110011111111: color_data = 12'b000001101111;
20'b01100111110100000000: color_data = 12'b000001101111;
20'b01100111110100000001: color_data = 12'b000001101111;
20'b01100111110100000010: color_data = 12'b000001101111;
20'b01100111110100000011: color_data = 12'b000001101111;
20'b01100111110100000100: color_data = 12'b000001101111;
20'b01100111110100000101: color_data = 12'b000001101111;
20'b01100111110100000110: color_data = 12'b000001101111;
20'b01100111110100000111: color_data = 12'b000001101111;
20'b01100111110100001000: color_data = 12'b000001101111;
20'b01100111110100001001: color_data = 12'b000001101111;
20'b01100111110100001010: color_data = 12'b000001101111;
20'b01100111110100001011: color_data = 12'b000001101111;
20'b01100111110100001111: color_data = 12'b000001101111;
20'b01100111110100010000: color_data = 12'b000001101111;
20'b01100111110100010001: color_data = 12'b000001101111;
20'b01100111110100010010: color_data = 12'b000001101111;
20'b01100111110100010011: color_data = 12'b000001101111;
20'b01100111110100010100: color_data = 12'b000001101111;
20'b01100111110100010101: color_data = 12'b000001101111;
20'b01100111110100010110: color_data = 12'b000001101111;
20'b01100111110100010111: color_data = 12'b000001101111;
20'b01100111110100011000: color_data = 12'b000001101111;
20'b01100111110100011001: color_data = 12'b000001101111;
20'b01100111110100011010: color_data = 12'b000001101111;
20'b01100111110100011011: color_data = 12'b000001101111;
20'b01100111110100011100: color_data = 12'b000001101111;
20'b01100111110100011101: color_data = 12'b000001101111;
20'b01100111110100011110: color_data = 12'b000001101111;
20'b01100111110100011111: color_data = 12'b000001101111;
20'b01100111110100100000: color_data = 12'b000001101111;
20'b01100111110100100100: color_data = 12'b000001101111;
20'b01100111110100100101: color_data = 12'b000001101111;
20'b01100111110100100110: color_data = 12'b000001101111;
20'b01100111110100100111: color_data = 12'b000001101111;
20'b01100111110100101000: color_data = 12'b000001101111;
20'b01100111110100101001: color_data = 12'b000001101111;
20'b01100111110100101010: color_data = 12'b000001101111;
20'b01100111110100101011: color_data = 12'b000001101111;
20'b01100111110100101100: color_data = 12'b000001101111;
20'b01100111110100101101: color_data = 12'b000001101111;
20'b01100111110100101110: color_data = 12'b000001101111;
20'b01100111110100101111: color_data = 12'b000001101111;
20'b01100111110100110000: color_data = 12'b000001101111;
20'b01100111110100110001: color_data = 12'b000001101111;
20'b01100111110100110010: color_data = 12'b000001101111;
20'b01100111110100110011: color_data = 12'b000001101111;
20'b01100111110100110100: color_data = 12'b000001101111;
20'b01100111110100110101: color_data = 12'b000001101111;
20'b01100111110100111001: color_data = 12'b000011110000;
20'b01100111110100111010: color_data = 12'b000011110000;
20'b01100111110100111011: color_data = 12'b000011110000;
20'b01100111110100111100: color_data = 12'b000011110000;
20'b01100111110100111101: color_data = 12'b000011110000;
20'b01100111110100111110: color_data = 12'b000011110000;
20'b01100111110100111111: color_data = 12'b000011110000;
20'b01100111110101000000: color_data = 12'b000011110000;
20'b01100111110101000001: color_data = 12'b000011110000;
20'b01100111110101000010: color_data = 12'b000011110000;
20'b01100111110101000011: color_data = 12'b000011110000;
20'b01100111110101000100: color_data = 12'b000011110000;
20'b01100111110101000101: color_data = 12'b000011110000;
20'b01100111110101000110: color_data = 12'b000011110000;
20'b01100111110101000111: color_data = 12'b000011110000;
20'b01100111110101001000: color_data = 12'b000011110000;
20'b01100111110101001001: color_data = 12'b000011110000;
20'b01100111110101001010: color_data = 12'b000011110000;
20'b01100111110101001110: color_data = 12'b000011110000;
20'b01100111110101001111: color_data = 12'b000011110000;
20'b01100111110101010000: color_data = 12'b000011110000;
20'b01100111110101010001: color_data = 12'b000011110000;
20'b01100111110101010010: color_data = 12'b000011110000;
20'b01100111110101010011: color_data = 12'b000011110000;
20'b01100111110101010100: color_data = 12'b000011110000;
20'b01100111110101010101: color_data = 12'b000011110000;
20'b01100111110101010110: color_data = 12'b000011110000;
20'b01100111110101010111: color_data = 12'b000011110000;
20'b01100111110101011000: color_data = 12'b000011110000;
20'b01100111110101011001: color_data = 12'b000011110000;
20'b01100111110101011010: color_data = 12'b000011110000;
20'b01100111110101011011: color_data = 12'b000011110000;
20'b01100111110101011100: color_data = 12'b000011110000;
20'b01100111110101011101: color_data = 12'b000011110000;
20'b01100111110101011110: color_data = 12'b000011110000;
20'b01100111110101011111: color_data = 12'b000011110000;
20'b01100111110101100011: color_data = 12'b111100001111;
20'b01100111110101100100: color_data = 12'b111100001111;
20'b01100111110101100101: color_data = 12'b111100001111;
20'b01100111110101100110: color_data = 12'b111100001111;
20'b01100111110101100111: color_data = 12'b111100001111;
20'b01100111110101101000: color_data = 12'b111100001111;
20'b01100111110101101001: color_data = 12'b111100001111;
20'b01100111110101101010: color_data = 12'b111100001111;
20'b01100111110101101011: color_data = 12'b111100001111;
20'b01100111110101101100: color_data = 12'b111100001111;
20'b01100111110101101101: color_data = 12'b111100001111;
20'b01100111110101101110: color_data = 12'b111100001111;
20'b01100111110101101111: color_data = 12'b111100001111;
20'b01100111110101110000: color_data = 12'b111100001111;
20'b01100111110101110001: color_data = 12'b111100001111;
20'b01100111110101110010: color_data = 12'b111100001111;
20'b01100111110101110011: color_data = 12'b111100001111;
20'b01100111110101110100: color_data = 12'b111100001111;
20'b01100111110101111000: color_data = 12'b111100001111;
20'b01100111110101111001: color_data = 12'b111100001111;
20'b01100111110101111010: color_data = 12'b111100001111;
20'b01100111110101111011: color_data = 12'b111100001111;
20'b01100111110101111100: color_data = 12'b111100001111;
20'b01100111110101111101: color_data = 12'b111100001111;
20'b01100111110101111110: color_data = 12'b111100001111;
20'b01100111110101111111: color_data = 12'b111100001111;
20'b01100111110110000000: color_data = 12'b111100001111;
20'b01100111110110000001: color_data = 12'b111100001111;
20'b01100111110110000010: color_data = 12'b111100001111;
20'b01100111110110000011: color_data = 12'b111100001111;
20'b01100111110110000100: color_data = 12'b111100001111;
20'b01100111110110000101: color_data = 12'b111100001111;
20'b01100111110110000110: color_data = 12'b111100001111;
20'b01100111110110000111: color_data = 12'b111100001111;
20'b01100111110110001000: color_data = 12'b111100001111;
20'b01100111110110001001: color_data = 12'b111100001111;
20'b01100111110110001101: color_data = 12'b111100000000;
20'b01100111110110001110: color_data = 12'b111100000000;
20'b01100111110110001111: color_data = 12'b111100000000;
20'b01100111110110010000: color_data = 12'b111100000000;
20'b01100111110110010001: color_data = 12'b111100000000;
20'b01100111110110010010: color_data = 12'b111100000000;
20'b01100111110110010011: color_data = 12'b111100000000;
20'b01100111110110010100: color_data = 12'b111100000000;
20'b01100111110110010101: color_data = 12'b111100000000;
20'b01100111110110010110: color_data = 12'b111100000000;
20'b01100111110110010111: color_data = 12'b111100000000;
20'b01100111110110011000: color_data = 12'b111100000000;
20'b01100111110110011001: color_data = 12'b111100000000;
20'b01100111110110011010: color_data = 12'b111100000000;
20'b01100111110110011011: color_data = 12'b111100000000;
20'b01100111110110011100: color_data = 12'b111100000000;
20'b01100111110110011101: color_data = 12'b111100000000;
20'b01100111110110011110: color_data = 12'b111100000000;
20'b01101000000011111010: color_data = 12'b000001101111;
20'b01101000000011111011: color_data = 12'b000001101111;
20'b01101000000011111100: color_data = 12'b000001101111;
20'b01101000000011111101: color_data = 12'b000001101111;
20'b01101000000011111110: color_data = 12'b000001101111;
20'b01101000000011111111: color_data = 12'b000001101111;
20'b01101000000100000000: color_data = 12'b000001101111;
20'b01101000000100000001: color_data = 12'b000001101111;
20'b01101000000100000010: color_data = 12'b000001101111;
20'b01101000000100000011: color_data = 12'b000001101111;
20'b01101000000100000100: color_data = 12'b000001101111;
20'b01101000000100000101: color_data = 12'b000001101111;
20'b01101000000100000110: color_data = 12'b000001101111;
20'b01101000000100000111: color_data = 12'b000001101111;
20'b01101000000100001000: color_data = 12'b000001101111;
20'b01101000000100001001: color_data = 12'b000001101111;
20'b01101000000100001010: color_data = 12'b000001101111;
20'b01101000000100001011: color_data = 12'b000001101111;
20'b01101000000100001111: color_data = 12'b000001101111;
20'b01101000000100010000: color_data = 12'b000001101111;
20'b01101000000100010001: color_data = 12'b000001101111;
20'b01101000000100010010: color_data = 12'b000001101111;
20'b01101000000100010011: color_data = 12'b000001101111;
20'b01101000000100010100: color_data = 12'b000001101111;
20'b01101000000100010101: color_data = 12'b000001101111;
20'b01101000000100010110: color_data = 12'b000001101111;
20'b01101000000100010111: color_data = 12'b000001101111;
20'b01101000000100011000: color_data = 12'b000001101111;
20'b01101000000100011001: color_data = 12'b000001101111;
20'b01101000000100011010: color_data = 12'b000001101111;
20'b01101000000100011011: color_data = 12'b000001101111;
20'b01101000000100011100: color_data = 12'b000001101111;
20'b01101000000100011101: color_data = 12'b000001101111;
20'b01101000000100011110: color_data = 12'b000001101111;
20'b01101000000100011111: color_data = 12'b000001101111;
20'b01101000000100100000: color_data = 12'b000001101111;
20'b01101000000100100100: color_data = 12'b000001101111;
20'b01101000000100100101: color_data = 12'b000001101111;
20'b01101000000100100110: color_data = 12'b000001101111;
20'b01101000000100100111: color_data = 12'b000001101111;
20'b01101000000100101000: color_data = 12'b000001101111;
20'b01101000000100101001: color_data = 12'b000001101111;
20'b01101000000100101010: color_data = 12'b000001101111;
20'b01101000000100101011: color_data = 12'b000001101111;
20'b01101000000100101100: color_data = 12'b000001101111;
20'b01101000000100101101: color_data = 12'b000001101111;
20'b01101000000100101110: color_data = 12'b000001101111;
20'b01101000000100101111: color_data = 12'b000001101111;
20'b01101000000100110000: color_data = 12'b000001101111;
20'b01101000000100110001: color_data = 12'b000001101111;
20'b01101000000100110010: color_data = 12'b000001101111;
20'b01101000000100110011: color_data = 12'b000001101111;
20'b01101000000100110100: color_data = 12'b000001101111;
20'b01101000000100110101: color_data = 12'b000001101111;
20'b01101000000100111001: color_data = 12'b000011110000;
20'b01101000000100111010: color_data = 12'b000011110000;
20'b01101000000100111011: color_data = 12'b000011110000;
20'b01101000000100111100: color_data = 12'b000011110000;
20'b01101000000100111101: color_data = 12'b000011110000;
20'b01101000000100111110: color_data = 12'b000011110000;
20'b01101000000100111111: color_data = 12'b000011110000;
20'b01101000000101000000: color_data = 12'b000011110000;
20'b01101000000101000001: color_data = 12'b000011110000;
20'b01101000000101000010: color_data = 12'b000011110000;
20'b01101000000101000011: color_data = 12'b000011110000;
20'b01101000000101000100: color_data = 12'b000011110000;
20'b01101000000101000101: color_data = 12'b000011110000;
20'b01101000000101000110: color_data = 12'b000011110000;
20'b01101000000101000111: color_data = 12'b000011110000;
20'b01101000000101001000: color_data = 12'b000011110000;
20'b01101000000101001001: color_data = 12'b000011110000;
20'b01101000000101001010: color_data = 12'b000011110000;
20'b01101000000101001110: color_data = 12'b000011110000;
20'b01101000000101001111: color_data = 12'b000011110000;
20'b01101000000101010000: color_data = 12'b000011110000;
20'b01101000000101010001: color_data = 12'b000011110000;
20'b01101000000101010010: color_data = 12'b000011110000;
20'b01101000000101010011: color_data = 12'b000011110000;
20'b01101000000101010100: color_data = 12'b000011110000;
20'b01101000000101010101: color_data = 12'b000011110000;
20'b01101000000101010110: color_data = 12'b000011110000;
20'b01101000000101010111: color_data = 12'b000011110000;
20'b01101000000101011000: color_data = 12'b000011110000;
20'b01101000000101011001: color_data = 12'b000011110000;
20'b01101000000101011010: color_data = 12'b000011110000;
20'b01101000000101011011: color_data = 12'b000011110000;
20'b01101000000101011100: color_data = 12'b000011110000;
20'b01101000000101011101: color_data = 12'b000011110000;
20'b01101000000101011110: color_data = 12'b000011110000;
20'b01101000000101011111: color_data = 12'b000011110000;
20'b01101000000101100011: color_data = 12'b111100001111;
20'b01101000000101100100: color_data = 12'b111100001111;
20'b01101000000101100101: color_data = 12'b111100001111;
20'b01101000000101100110: color_data = 12'b111100001111;
20'b01101000000101100111: color_data = 12'b111100001111;
20'b01101000000101101000: color_data = 12'b111100001111;
20'b01101000000101101001: color_data = 12'b111100001111;
20'b01101000000101101010: color_data = 12'b111100001111;
20'b01101000000101101011: color_data = 12'b111100001111;
20'b01101000000101101100: color_data = 12'b111100001111;
20'b01101000000101101101: color_data = 12'b111100001111;
20'b01101000000101101110: color_data = 12'b111100001111;
20'b01101000000101101111: color_data = 12'b111100001111;
20'b01101000000101110000: color_data = 12'b111100001111;
20'b01101000000101110001: color_data = 12'b111100001111;
20'b01101000000101110010: color_data = 12'b111100001111;
20'b01101000000101110011: color_data = 12'b111100001111;
20'b01101000000101110100: color_data = 12'b111100001111;
20'b01101000000101111000: color_data = 12'b111100001111;
20'b01101000000101111001: color_data = 12'b111100001111;
20'b01101000000101111010: color_data = 12'b111100001111;
20'b01101000000101111011: color_data = 12'b111100001111;
20'b01101000000101111100: color_data = 12'b111100001111;
20'b01101000000101111101: color_data = 12'b111100001111;
20'b01101000000101111110: color_data = 12'b111100001111;
20'b01101000000101111111: color_data = 12'b111100001111;
20'b01101000000110000000: color_data = 12'b111100001111;
20'b01101000000110000001: color_data = 12'b111100001111;
20'b01101000000110000010: color_data = 12'b111100001111;
20'b01101000000110000011: color_data = 12'b111100001111;
20'b01101000000110000100: color_data = 12'b111100001111;
20'b01101000000110000101: color_data = 12'b111100001111;
20'b01101000000110000110: color_data = 12'b111100001111;
20'b01101000000110000111: color_data = 12'b111100001111;
20'b01101000000110001000: color_data = 12'b111100001111;
20'b01101000000110001001: color_data = 12'b111100001111;
20'b01101000000110001101: color_data = 12'b111100000000;
20'b01101000000110001110: color_data = 12'b111100000000;
20'b01101000000110001111: color_data = 12'b111100000000;
20'b01101000000110010000: color_data = 12'b111100000000;
20'b01101000000110010001: color_data = 12'b111100000000;
20'b01101000000110010010: color_data = 12'b111100000000;
20'b01101000000110010011: color_data = 12'b111100000000;
20'b01101000000110010100: color_data = 12'b111100000000;
20'b01101000000110010101: color_data = 12'b111100000000;
20'b01101000000110010110: color_data = 12'b111100000000;
20'b01101000000110010111: color_data = 12'b111100000000;
20'b01101000000110011000: color_data = 12'b111100000000;
20'b01101000000110011001: color_data = 12'b111100000000;
20'b01101000000110011010: color_data = 12'b111100000000;
20'b01101000000110011011: color_data = 12'b111100000000;
20'b01101000000110011100: color_data = 12'b111100000000;
20'b01101000000110011101: color_data = 12'b111100000000;
20'b01101000000110011110: color_data = 12'b111100000000;
20'b01101000010011111010: color_data = 12'b000001101111;
20'b01101000010011111011: color_data = 12'b000001101111;
20'b01101000010011111100: color_data = 12'b000001101111;
20'b01101000010011111101: color_data = 12'b000001101111;
20'b01101000010011111110: color_data = 12'b000001101111;
20'b01101000010011111111: color_data = 12'b000001101111;
20'b01101000010100000000: color_data = 12'b000001101111;
20'b01101000010100000001: color_data = 12'b000001101111;
20'b01101000010100000010: color_data = 12'b000001101111;
20'b01101000010100000011: color_data = 12'b000001101111;
20'b01101000010100000100: color_data = 12'b000001101111;
20'b01101000010100000101: color_data = 12'b000001101111;
20'b01101000010100000110: color_data = 12'b000001101111;
20'b01101000010100000111: color_data = 12'b000001101111;
20'b01101000010100001000: color_data = 12'b000001101111;
20'b01101000010100001001: color_data = 12'b000001101111;
20'b01101000010100001010: color_data = 12'b000001101111;
20'b01101000010100001011: color_data = 12'b000001101111;
20'b01101000010100001111: color_data = 12'b000001101111;
20'b01101000010100010000: color_data = 12'b000001101111;
20'b01101000010100010001: color_data = 12'b000001101111;
20'b01101000010100010010: color_data = 12'b000001101111;
20'b01101000010100010011: color_data = 12'b000001101111;
20'b01101000010100010100: color_data = 12'b000001101111;
20'b01101000010100010101: color_data = 12'b000001101111;
20'b01101000010100010110: color_data = 12'b000001101111;
20'b01101000010100010111: color_data = 12'b000001101111;
20'b01101000010100011000: color_data = 12'b000001101111;
20'b01101000010100011001: color_data = 12'b000001101111;
20'b01101000010100011010: color_data = 12'b000001101111;
20'b01101000010100011011: color_data = 12'b000001101111;
20'b01101000010100011100: color_data = 12'b000001101111;
20'b01101000010100011101: color_data = 12'b000001101111;
20'b01101000010100011110: color_data = 12'b000001101111;
20'b01101000010100011111: color_data = 12'b000001101111;
20'b01101000010100100000: color_data = 12'b000001101111;
20'b01101000010100100100: color_data = 12'b000001101111;
20'b01101000010100100101: color_data = 12'b000001101111;
20'b01101000010100100110: color_data = 12'b000001101111;
20'b01101000010100100111: color_data = 12'b000001101111;
20'b01101000010100101000: color_data = 12'b000001101111;
20'b01101000010100101001: color_data = 12'b000001101111;
20'b01101000010100101010: color_data = 12'b000001101111;
20'b01101000010100101011: color_data = 12'b000001101111;
20'b01101000010100101100: color_data = 12'b000001101111;
20'b01101000010100101101: color_data = 12'b000001101111;
20'b01101000010100101110: color_data = 12'b000001101111;
20'b01101000010100101111: color_data = 12'b000001101111;
20'b01101000010100110000: color_data = 12'b000001101111;
20'b01101000010100110001: color_data = 12'b000001101111;
20'b01101000010100110010: color_data = 12'b000001101111;
20'b01101000010100110011: color_data = 12'b000001101111;
20'b01101000010100110100: color_data = 12'b000001101111;
20'b01101000010100110101: color_data = 12'b000001101111;
20'b01101000010100111001: color_data = 12'b000011110000;
20'b01101000010100111010: color_data = 12'b000011110000;
20'b01101000010100111011: color_data = 12'b000011110000;
20'b01101000010100111100: color_data = 12'b000011110000;
20'b01101000010100111101: color_data = 12'b000011110000;
20'b01101000010100111110: color_data = 12'b000011110000;
20'b01101000010100111111: color_data = 12'b000011110000;
20'b01101000010101000000: color_data = 12'b000011110000;
20'b01101000010101000001: color_data = 12'b000011110000;
20'b01101000010101000010: color_data = 12'b000011110000;
20'b01101000010101000011: color_data = 12'b000011110000;
20'b01101000010101000100: color_data = 12'b000011110000;
20'b01101000010101000101: color_data = 12'b000011110000;
20'b01101000010101000110: color_data = 12'b000011110000;
20'b01101000010101000111: color_data = 12'b000011110000;
20'b01101000010101001000: color_data = 12'b000011110000;
20'b01101000010101001001: color_data = 12'b000011110000;
20'b01101000010101001010: color_data = 12'b000011110000;
20'b01101000010101001110: color_data = 12'b000011110000;
20'b01101000010101001111: color_data = 12'b000011110000;
20'b01101000010101010000: color_data = 12'b000011110000;
20'b01101000010101010001: color_data = 12'b000011110000;
20'b01101000010101010010: color_data = 12'b000011110000;
20'b01101000010101010011: color_data = 12'b000011110000;
20'b01101000010101010100: color_data = 12'b000011110000;
20'b01101000010101010101: color_data = 12'b000011110000;
20'b01101000010101010110: color_data = 12'b000011110000;
20'b01101000010101010111: color_data = 12'b000011110000;
20'b01101000010101011000: color_data = 12'b000011110000;
20'b01101000010101011001: color_data = 12'b000011110000;
20'b01101000010101011010: color_data = 12'b000011110000;
20'b01101000010101011011: color_data = 12'b000011110000;
20'b01101000010101011100: color_data = 12'b000011110000;
20'b01101000010101011101: color_data = 12'b000011110000;
20'b01101000010101011110: color_data = 12'b000011110000;
20'b01101000010101011111: color_data = 12'b000011110000;
20'b01101000010101100011: color_data = 12'b111100001111;
20'b01101000010101100100: color_data = 12'b111100001111;
20'b01101000010101100101: color_data = 12'b111100001111;
20'b01101000010101100110: color_data = 12'b111100001111;
20'b01101000010101100111: color_data = 12'b111100001111;
20'b01101000010101101000: color_data = 12'b111100001111;
20'b01101000010101101001: color_data = 12'b111100001111;
20'b01101000010101101010: color_data = 12'b111100001111;
20'b01101000010101101011: color_data = 12'b111100001111;
20'b01101000010101101100: color_data = 12'b111100001111;
20'b01101000010101101101: color_data = 12'b111100001111;
20'b01101000010101101110: color_data = 12'b111100001111;
20'b01101000010101101111: color_data = 12'b111100001111;
20'b01101000010101110000: color_data = 12'b111100001111;
20'b01101000010101110001: color_data = 12'b111100001111;
20'b01101000010101110010: color_data = 12'b111100001111;
20'b01101000010101110011: color_data = 12'b111100001111;
20'b01101000010101110100: color_data = 12'b111100001111;
20'b01101000010101111000: color_data = 12'b111100001111;
20'b01101000010101111001: color_data = 12'b111100001111;
20'b01101000010101111010: color_data = 12'b111100001111;
20'b01101000010101111011: color_data = 12'b111100001111;
20'b01101000010101111100: color_data = 12'b111100001111;
20'b01101000010101111101: color_data = 12'b111100001111;
20'b01101000010101111110: color_data = 12'b111100001111;
20'b01101000010101111111: color_data = 12'b111100001111;
20'b01101000010110000000: color_data = 12'b111100001111;
20'b01101000010110000001: color_data = 12'b111100001111;
20'b01101000010110000010: color_data = 12'b111100001111;
20'b01101000010110000011: color_data = 12'b111100001111;
20'b01101000010110000100: color_data = 12'b111100001111;
20'b01101000010110000101: color_data = 12'b111100001111;
20'b01101000010110000110: color_data = 12'b111100001111;
20'b01101000010110000111: color_data = 12'b111100001111;
20'b01101000010110001000: color_data = 12'b111100001111;
20'b01101000010110001001: color_data = 12'b111100001111;
20'b01101000010110001101: color_data = 12'b111100000000;
20'b01101000010110001110: color_data = 12'b111100000000;
20'b01101000010110001111: color_data = 12'b111100000000;
20'b01101000010110010000: color_data = 12'b111100000000;
20'b01101000010110010001: color_data = 12'b111100000000;
20'b01101000010110010010: color_data = 12'b111100000000;
20'b01101000010110010011: color_data = 12'b111100000000;
20'b01101000010110010100: color_data = 12'b111100000000;
20'b01101000010110010101: color_data = 12'b111100000000;
20'b01101000010110010110: color_data = 12'b111100000000;
20'b01101000010110010111: color_data = 12'b111100000000;
20'b01101000010110011000: color_data = 12'b111100000000;
20'b01101000010110011001: color_data = 12'b111100000000;
20'b01101000010110011010: color_data = 12'b111100000000;
20'b01101000010110011011: color_data = 12'b111100000000;
20'b01101000010110011100: color_data = 12'b111100000000;
20'b01101000010110011101: color_data = 12'b111100000000;
20'b01101000010110011110: color_data = 12'b111100000000;
20'b01101001010011111010: color_data = 12'b111101110000;
20'b01101001010011111011: color_data = 12'b111101110000;
20'b01101001010011111100: color_data = 12'b111101110000;
20'b01101001010011111101: color_data = 12'b111101110000;
20'b01101001010011111110: color_data = 12'b111101110000;
20'b01101001010011111111: color_data = 12'b111101110000;
20'b01101001010100000000: color_data = 12'b111101110000;
20'b01101001010100000001: color_data = 12'b111101110000;
20'b01101001010100000010: color_data = 12'b111101110000;
20'b01101001010100000011: color_data = 12'b111101110000;
20'b01101001010100000100: color_data = 12'b111101110000;
20'b01101001010100000101: color_data = 12'b111101110000;
20'b01101001010100000110: color_data = 12'b111101110000;
20'b01101001010100000111: color_data = 12'b111101110000;
20'b01101001010100001000: color_data = 12'b111101110000;
20'b01101001010100001001: color_data = 12'b111101110000;
20'b01101001010100001010: color_data = 12'b111101110000;
20'b01101001010100001011: color_data = 12'b111101110000;
20'b01101001010100001111: color_data = 12'b111101110000;
20'b01101001010100010000: color_data = 12'b111101110000;
20'b01101001010100010001: color_data = 12'b111101110000;
20'b01101001010100010010: color_data = 12'b111101110000;
20'b01101001010100010011: color_data = 12'b111101110000;
20'b01101001010100010100: color_data = 12'b111101110000;
20'b01101001010100010101: color_data = 12'b111101110000;
20'b01101001010100010110: color_data = 12'b111101110000;
20'b01101001010100010111: color_data = 12'b111101110000;
20'b01101001010100011000: color_data = 12'b111101110000;
20'b01101001010100011001: color_data = 12'b111101110000;
20'b01101001010100011010: color_data = 12'b111101110000;
20'b01101001010100011011: color_data = 12'b111101110000;
20'b01101001010100011100: color_data = 12'b111101110000;
20'b01101001010100011101: color_data = 12'b111101110000;
20'b01101001010100011110: color_data = 12'b111101110000;
20'b01101001010100011111: color_data = 12'b111101110000;
20'b01101001010100100000: color_data = 12'b111101110000;
20'b01101001010100100100: color_data = 12'b111101110000;
20'b01101001010100100101: color_data = 12'b111101110000;
20'b01101001010100100110: color_data = 12'b111101110000;
20'b01101001010100100111: color_data = 12'b111101110000;
20'b01101001010100101000: color_data = 12'b111101110000;
20'b01101001010100101001: color_data = 12'b111101110000;
20'b01101001010100101010: color_data = 12'b111101110000;
20'b01101001010100101011: color_data = 12'b111101110000;
20'b01101001010100101100: color_data = 12'b111101110000;
20'b01101001010100101101: color_data = 12'b111101110000;
20'b01101001010100101110: color_data = 12'b111101110000;
20'b01101001010100101111: color_data = 12'b111101110000;
20'b01101001010100110000: color_data = 12'b111101110000;
20'b01101001010100110001: color_data = 12'b111101110000;
20'b01101001010100110010: color_data = 12'b111101110000;
20'b01101001010100110011: color_data = 12'b111101110000;
20'b01101001010100110100: color_data = 12'b111101110000;
20'b01101001010100110101: color_data = 12'b111101110000;
20'b01101001010100111001: color_data = 12'b111101110000;
20'b01101001010100111010: color_data = 12'b111101110000;
20'b01101001010100111011: color_data = 12'b111101110000;
20'b01101001010100111100: color_data = 12'b111101110000;
20'b01101001010100111101: color_data = 12'b111101110000;
20'b01101001010100111110: color_data = 12'b111101110000;
20'b01101001010100111111: color_data = 12'b111101110000;
20'b01101001010101000000: color_data = 12'b111101110000;
20'b01101001010101000001: color_data = 12'b111101110000;
20'b01101001010101000010: color_data = 12'b111101110000;
20'b01101001010101000011: color_data = 12'b111101110000;
20'b01101001010101000100: color_data = 12'b111101110000;
20'b01101001010101000101: color_data = 12'b111101110000;
20'b01101001010101000110: color_data = 12'b111101110000;
20'b01101001010101000111: color_data = 12'b111101110000;
20'b01101001010101001000: color_data = 12'b111101110000;
20'b01101001010101001001: color_data = 12'b111101110000;
20'b01101001010101001010: color_data = 12'b111101110000;
20'b01101001010101001110: color_data = 12'b000011110000;
20'b01101001010101001111: color_data = 12'b000011110000;
20'b01101001010101010000: color_data = 12'b000011110000;
20'b01101001010101010001: color_data = 12'b000011110000;
20'b01101001010101010010: color_data = 12'b000011110000;
20'b01101001010101010011: color_data = 12'b000011110000;
20'b01101001010101010100: color_data = 12'b000011110000;
20'b01101001010101010101: color_data = 12'b000011110000;
20'b01101001010101010110: color_data = 12'b000011110000;
20'b01101001010101010111: color_data = 12'b000011110000;
20'b01101001010101011000: color_data = 12'b000011110000;
20'b01101001010101011001: color_data = 12'b000011110000;
20'b01101001010101011010: color_data = 12'b000011110000;
20'b01101001010101011011: color_data = 12'b000011110000;
20'b01101001010101011100: color_data = 12'b000011110000;
20'b01101001010101011101: color_data = 12'b000011110000;
20'b01101001010101011110: color_data = 12'b000011110000;
20'b01101001010101011111: color_data = 12'b000011110000;
20'b01101001010101100011: color_data = 12'b111100001111;
20'b01101001010101100100: color_data = 12'b111100001111;
20'b01101001010101100101: color_data = 12'b111100001111;
20'b01101001010101100110: color_data = 12'b111100001111;
20'b01101001010101100111: color_data = 12'b111100001111;
20'b01101001010101101000: color_data = 12'b111100001111;
20'b01101001010101101001: color_data = 12'b111100001111;
20'b01101001010101101010: color_data = 12'b111100001111;
20'b01101001010101101011: color_data = 12'b111100001111;
20'b01101001010101101100: color_data = 12'b111100001111;
20'b01101001010101101101: color_data = 12'b111100001111;
20'b01101001010101101110: color_data = 12'b111100001111;
20'b01101001010101101111: color_data = 12'b111100001111;
20'b01101001010101110000: color_data = 12'b111100001111;
20'b01101001010101110001: color_data = 12'b111100001111;
20'b01101001010101110010: color_data = 12'b111100001111;
20'b01101001010101110011: color_data = 12'b111100001111;
20'b01101001010101110100: color_data = 12'b111100001111;
20'b01101001010101111000: color_data = 12'b111100000000;
20'b01101001010101111001: color_data = 12'b111100000000;
20'b01101001010101111010: color_data = 12'b111100000000;
20'b01101001010101111011: color_data = 12'b111100000000;
20'b01101001010101111100: color_data = 12'b111100000000;
20'b01101001010101111101: color_data = 12'b111100000000;
20'b01101001010101111110: color_data = 12'b111100000000;
20'b01101001010101111111: color_data = 12'b111100000000;
20'b01101001010110000000: color_data = 12'b111100000000;
20'b01101001010110000001: color_data = 12'b111100000000;
20'b01101001010110000010: color_data = 12'b111100000000;
20'b01101001010110000011: color_data = 12'b111100000000;
20'b01101001010110000100: color_data = 12'b111100000000;
20'b01101001010110000101: color_data = 12'b111100000000;
20'b01101001010110000110: color_data = 12'b111100000000;
20'b01101001010110000111: color_data = 12'b111100000000;
20'b01101001010110001000: color_data = 12'b111100000000;
20'b01101001010110001001: color_data = 12'b111100000000;
20'b01101001010110001101: color_data = 12'b111100000000;
20'b01101001010110001110: color_data = 12'b111100000000;
20'b01101001010110001111: color_data = 12'b111100000000;
20'b01101001010110010000: color_data = 12'b111100000000;
20'b01101001010110010001: color_data = 12'b111100000000;
20'b01101001010110010010: color_data = 12'b111100000000;
20'b01101001010110010011: color_data = 12'b111100000000;
20'b01101001010110010100: color_data = 12'b111100000000;
20'b01101001010110010101: color_data = 12'b111100000000;
20'b01101001010110010110: color_data = 12'b111100000000;
20'b01101001010110010111: color_data = 12'b111100000000;
20'b01101001010110011000: color_data = 12'b111100000000;
20'b01101001010110011001: color_data = 12'b111100000000;
20'b01101001010110011010: color_data = 12'b111100000000;
20'b01101001010110011011: color_data = 12'b111100000000;
20'b01101001010110011100: color_data = 12'b111100000000;
20'b01101001010110011101: color_data = 12'b111100000000;
20'b01101001010110011110: color_data = 12'b111100000000;
20'b01101001100011111010: color_data = 12'b111101110000;
20'b01101001100011111011: color_data = 12'b111101110000;
20'b01101001100011111100: color_data = 12'b111101110000;
20'b01101001100011111101: color_data = 12'b111101110000;
20'b01101001100011111110: color_data = 12'b111101110000;
20'b01101001100011111111: color_data = 12'b111101110000;
20'b01101001100100000000: color_data = 12'b111101110000;
20'b01101001100100000001: color_data = 12'b111101110000;
20'b01101001100100000010: color_data = 12'b111101110000;
20'b01101001100100000011: color_data = 12'b111101110000;
20'b01101001100100000100: color_data = 12'b111101110000;
20'b01101001100100000101: color_data = 12'b111101110000;
20'b01101001100100000110: color_data = 12'b111101110000;
20'b01101001100100000111: color_data = 12'b111101110000;
20'b01101001100100001000: color_data = 12'b111101110000;
20'b01101001100100001001: color_data = 12'b111101110000;
20'b01101001100100001010: color_data = 12'b111101110000;
20'b01101001100100001011: color_data = 12'b111101110000;
20'b01101001100100001111: color_data = 12'b111101110000;
20'b01101001100100010000: color_data = 12'b111101110000;
20'b01101001100100010001: color_data = 12'b111101110000;
20'b01101001100100010010: color_data = 12'b111101110000;
20'b01101001100100010011: color_data = 12'b111101110000;
20'b01101001100100010100: color_data = 12'b111101110000;
20'b01101001100100010101: color_data = 12'b111101110000;
20'b01101001100100010110: color_data = 12'b111101110000;
20'b01101001100100010111: color_data = 12'b111101110000;
20'b01101001100100011000: color_data = 12'b111101110000;
20'b01101001100100011001: color_data = 12'b111101110000;
20'b01101001100100011010: color_data = 12'b111101110000;
20'b01101001100100011011: color_data = 12'b111101110000;
20'b01101001100100011100: color_data = 12'b111101110000;
20'b01101001100100011101: color_data = 12'b111101110000;
20'b01101001100100011110: color_data = 12'b111101110000;
20'b01101001100100011111: color_data = 12'b111101110000;
20'b01101001100100100000: color_data = 12'b111101110000;
20'b01101001100100100100: color_data = 12'b111101110000;
20'b01101001100100100101: color_data = 12'b111101110000;
20'b01101001100100100110: color_data = 12'b111101110000;
20'b01101001100100100111: color_data = 12'b111101110000;
20'b01101001100100101000: color_data = 12'b111101110000;
20'b01101001100100101001: color_data = 12'b111101110000;
20'b01101001100100101010: color_data = 12'b111101110000;
20'b01101001100100101011: color_data = 12'b111101110000;
20'b01101001100100101100: color_data = 12'b111101110000;
20'b01101001100100101101: color_data = 12'b111101110000;
20'b01101001100100101110: color_data = 12'b111101110000;
20'b01101001100100101111: color_data = 12'b111101110000;
20'b01101001100100110000: color_data = 12'b111101110000;
20'b01101001100100110001: color_data = 12'b111101110000;
20'b01101001100100110010: color_data = 12'b111101110000;
20'b01101001100100110011: color_data = 12'b111101110000;
20'b01101001100100110100: color_data = 12'b111101110000;
20'b01101001100100110101: color_data = 12'b111101110000;
20'b01101001100100111001: color_data = 12'b111101110000;
20'b01101001100100111010: color_data = 12'b111101110000;
20'b01101001100100111011: color_data = 12'b111101110000;
20'b01101001100100111100: color_data = 12'b111101110000;
20'b01101001100100111101: color_data = 12'b111101110000;
20'b01101001100100111110: color_data = 12'b111101110000;
20'b01101001100100111111: color_data = 12'b111101110000;
20'b01101001100101000000: color_data = 12'b111101110000;
20'b01101001100101000001: color_data = 12'b111101110000;
20'b01101001100101000010: color_data = 12'b111101110000;
20'b01101001100101000011: color_data = 12'b111101110000;
20'b01101001100101000100: color_data = 12'b111101110000;
20'b01101001100101000101: color_data = 12'b111101110000;
20'b01101001100101000110: color_data = 12'b111101110000;
20'b01101001100101000111: color_data = 12'b111101110000;
20'b01101001100101001000: color_data = 12'b111101110000;
20'b01101001100101001001: color_data = 12'b111101110000;
20'b01101001100101001010: color_data = 12'b111101110000;
20'b01101001100101001110: color_data = 12'b000011110000;
20'b01101001100101001111: color_data = 12'b000011110000;
20'b01101001100101010000: color_data = 12'b000011110000;
20'b01101001100101010001: color_data = 12'b000011110000;
20'b01101001100101010010: color_data = 12'b000011110000;
20'b01101001100101010011: color_data = 12'b000011110000;
20'b01101001100101010100: color_data = 12'b000011110000;
20'b01101001100101010101: color_data = 12'b000011110000;
20'b01101001100101010110: color_data = 12'b000011110000;
20'b01101001100101010111: color_data = 12'b000011110000;
20'b01101001100101011000: color_data = 12'b000011110000;
20'b01101001100101011001: color_data = 12'b000011110000;
20'b01101001100101011010: color_data = 12'b000011110000;
20'b01101001100101011011: color_data = 12'b000011110000;
20'b01101001100101011100: color_data = 12'b000011110000;
20'b01101001100101011101: color_data = 12'b000011110000;
20'b01101001100101011110: color_data = 12'b000011110000;
20'b01101001100101011111: color_data = 12'b000011110000;
20'b01101001100101100011: color_data = 12'b111100001111;
20'b01101001100101100100: color_data = 12'b111100001111;
20'b01101001100101100101: color_data = 12'b111100001111;
20'b01101001100101100110: color_data = 12'b111100001111;
20'b01101001100101100111: color_data = 12'b111100001111;
20'b01101001100101101000: color_data = 12'b111100001111;
20'b01101001100101101001: color_data = 12'b111100001111;
20'b01101001100101101010: color_data = 12'b111100001111;
20'b01101001100101101011: color_data = 12'b111100001111;
20'b01101001100101101100: color_data = 12'b111100001111;
20'b01101001100101101101: color_data = 12'b111100001111;
20'b01101001100101101110: color_data = 12'b111100001111;
20'b01101001100101101111: color_data = 12'b111100001111;
20'b01101001100101110000: color_data = 12'b111100001111;
20'b01101001100101110001: color_data = 12'b111100001111;
20'b01101001100101110010: color_data = 12'b111100001111;
20'b01101001100101110011: color_data = 12'b111100001111;
20'b01101001100101110100: color_data = 12'b111100001111;
20'b01101001100101111000: color_data = 12'b111100000000;
20'b01101001100101111001: color_data = 12'b111100000000;
20'b01101001100101111010: color_data = 12'b111100000000;
20'b01101001100101111011: color_data = 12'b111100000000;
20'b01101001100101111100: color_data = 12'b111100000000;
20'b01101001100101111101: color_data = 12'b111100000000;
20'b01101001100101111110: color_data = 12'b111100000000;
20'b01101001100101111111: color_data = 12'b111100000000;
20'b01101001100110000000: color_data = 12'b111100000000;
20'b01101001100110000001: color_data = 12'b111100000000;
20'b01101001100110000010: color_data = 12'b111100000000;
20'b01101001100110000011: color_data = 12'b111100000000;
20'b01101001100110000100: color_data = 12'b111100000000;
20'b01101001100110000101: color_data = 12'b111100000000;
20'b01101001100110000110: color_data = 12'b111100000000;
20'b01101001100110000111: color_data = 12'b111100000000;
20'b01101001100110001000: color_data = 12'b111100000000;
20'b01101001100110001001: color_data = 12'b111100000000;
20'b01101001100110001101: color_data = 12'b111100000000;
20'b01101001100110001110: color_data = 12'b111100000000;
20'b01101001100110001111: color_data = 12'b111100000000;
20'b01101001100110010000: color_data = 12'b111100000000;
20'b01101001100110010001: color_data = 12'b111100000000;
20'b01101001100110010010: color_data = 12'b111100000000;
20'b01101001100110010011: color_data = 12'b111100000000;
20'b01101001100110010100: color_data = 12'b111100000000;
20'b01101001100110010101: color_data = 12'b111100000000;
20'b01101001100110010110: color_data = 12'b111100000000;
20'b01101001100110010111: color_data = 12'b111100000000;
20'b01101001100110011000: color_data = 12'b111100000000;
20'b01101001100110011001: color_data = 12'b111100000000;
20'b01101001100110011010: color_data = 12'b111100000000;
20'b01101001100110011011: color_data = 12'b111100000000;
20'b01101001100110011100: color_data = 12'b111100000000;
20'b01101001100110011101: color_data = 12'b111100000000;
20'b01101001100110011110: color_data = 12'b111100000000;
20'b01101001110011111010: color_data = 12'b111101110000;
20'b01101001110011111011: color_data = 12'b111101110000;
20'b01101001110011111100: color_data = 12'b111101110000;
20'b01101001110011111101: color_data = 12'b111101110000;
20'b01101001110011111110: color_data = 12'b111101110000;
20'b01101001110011111111: color_data = 12'b111101110000;
20'b01101001110100000000: color_data = 12'b111101110000;
20'b01101001110100000001: color_data = 12'b111101110000;
20'b01101001110100000010: color_data = 12'b111101110000;
20'b01101001110100000011: color_data = 12'b111101110000;
20'b01101001110100000100: color_data = 12'b111101110000;
20'b01101001110100000101: color_data = 12'b111101110000;
20'b01101001110100000110: color_data = 12'b111101110000;
20'b01101001110100000111: color_data = 12'b111101110000;
20'b01101001110100001000: color_data = 12'b111101110000;
20'b01101001110100001001: color_data = 12'b111101110000;
20'b01101001110100001010: color_data = 12'b111101110000;
20'b01101001110100001011: color_data = 12'b111101110000;
20'b01101001110100001111: color_data = 12'b111101110000;
20'b01101001110100010000: color_data = 12'b111101110000;
20'b01101001110100010001: color_data = 12'b111101110000;
20'b01101001110100010010: color_data = 12'b111101110000;
20'b01101001110100010011: color_data = 12'b111101110000;
20'b01101001110100010100: color_data = 12'b111101110000;
20'b01101001110100010101: color_data = 12'b111101110000;
20'b01101001110100010110: color_data = 12'b111101110000;
20'b01101001110100010111: color_data = 12'b111101110000;
20'b01101001110100011000: color_data = 12'b111101110000;
20'b01101001110100011001: color_data = 12'b111101110000;
20'b01101001110100011010: color_data = 12'b111101110000;
20'b01101001110100011011: color_data = 12'b111101110000;
20'b01101001110100011100: color_data = 12'b111101110000;
20'b01101001110100011101: color_data = 12'b111101110000;
20'b01101001110100011110: color_data = 12'b111101110000;
20'b01101001110100011111: color_data = 12'b111101110000;
20'b01101001110100100000: color_data = 12'b111101110000;
20'b01101001110100100100: color_data = 12'b111101110000;
20'b01101001110100100101: color_data = 12'b111101110000;
20'b01101001110100100110: color_data = 12'b111101110000;
20'b01101001110100100111: color_data = 12'b111101110000;
20'b01101001110100101000: color_data = 12'b111101110000;
20'b01101001110100101001: color_data = 12'b111101110000;
20'b01101001110100101010: color_data = 12'b111101110000;
20'b01101001110100101011: color_data = 12'b111101110000;
20'b01101001110100101100: color_data = 12'b111101110000;
20'b01101001110100101101: color_data = 12'b111101110000;
20'b01101001110100101110: color_data = 12'b111101110000;
20'b01101001110100101111: color_data = 12'b111101110000;
20'b01101001110100110000: color_data = 12'b111101110000;
20'b01101001110100110001: color_data = 12'b111101110000;
20'b01101001110100110010: color_data = 12'b111101110000;
20'b01101001110100110011: color_data = 12'b111101110000;
20'b01101001110100110100: color_data = 12'b111101110000;
20'b01101001110100110101: color_data = 12'b111101110000;
20'b01101001110100111001: color_data = 12'b111101110000;
20'b01101001110100111010: color_data = 12'b111101110000;
20'b01101001110100111011: color_data = 12'b111101110000;
20'b01101001110100111100: color_data = 12'b111101110000;
20'b01101001110100111101: color_data = 12'b111101110000;
20'b01101001110100111110: color_data = 12'b111101110000;
20'b01101001110100111111: color_data = 12'b111101110000;
20'b01101001110101000000: color_data = 12'b111101110000;
20'b01101001110101000001: color_data = 12'b111101110000;
20'b01101001110101000010: color_data = 12'b111101110000;
20'b01101001110101000011: color_data = 12'b111101110000;
20'b01101001110101000100: color_data = 12'b111101110000;
20'b01101001110101000101: color_data = 12'b111101110000;
20'b01101001110101000110: color_data = 12'b111101110000;
20'b01101001110101000111: color_data = 12'b111101110000;
20'b01101001110101001000: color_data = 12'b111101110000;
20'b01101001110101001001: color_data = 12'b111101110000;
20'b01101001110101001010: color_data = 12'b111101110000;
20'b01101001110101001110: color_data = 12'b000011110000;
20'b01101001110101001111: color_data = 12'b000011110000;
20'b01101001110101010000: color_data = 12'b000011110000;
20'b01101001110101010001: color_data = 12'b000011110000;
20'b01101001110101010010: color_data = 12'b000011110000;
20'b01101001110101010011: color_data = 12'b000011110000;
20'b01101001110101010100: color_data = 12'b000011110000;
20'b01101001110101010101: color_data = 12'b000011110000;
20'b01101001110101010110: color_data = 12'b000011110000;
20'b01101001110101010111: color_data = 12'b000011110000;
20'b01101001110101011000: color_data = 12'b000011110000;
20'b01101001110101011001: color_data = 12'b000011110000;
20'b01101001110101011010: color_data = 12'b000011110000;
20'b01101001110101011011: color_data = 12'b000011110000;
20'b01101001110101011100: color_data = 12'b000011110000;
20'b01101001110101011101: color_data = 12'b000011110000;
20'b01101001110101011110: color_data = 12'b000011110000;
20'b01101001110101011111: color_data = 12'b000011110000;
20'b01101001110101100011: color_data = 12'b111100001111;
20'b01101001110101100100: color_data = 12'b111100001111;
20'b01101001110101100101: color_data = 12'b111100001111;
20'b01101001110101100110: color_data = 12'b111100001111;
20'b01101001110101100111: color_data = 12'b111100001111;
20'b01101001110101101000: color_data = 12'b111100001111;
20'b01101001110101101001: color_data = 12'b111100001111;
20'b01101001110101101010: color_data = 12'b111100001111;
20'b01101001110101101011: color_data = 12'b111100001111;
20'b01101001110101101100: color_data = 12'b111100001111;
20'b01101001110101101101: color_data = 12'b111100001111;
20'b01101001110101101110: color_data = 12'b111100001111;
20'b01101001110101101111: color_data = 12'b111100001111;
20'b01101001110101110000: color_data = 12'b111100001111;
20'b01101001110101110001: color_data = 12'b111100001111;
20'b01101001110101110010: color_data = 12'b111100001111;
20'b01101001110101110011: color_data = 12'b111100001111;
20'b01101001110101110100: color_data = 12'b111100001111;
20'b01101001110101111000: color_data = 12'b111100000000;
20'b01101001110101111001: color_data = 12'b111100000000;
20'b01101001110101111010: color_data = 12'b111100000000;
20'b01101001110101111011: color_data = 12'b111100000000;
20'b01101001110101111100: color_data = 12'b111100000000;
20'b01101001110101111101: color_data = 12'b111100000000;
20'b01101001110101111110: color_data = 12'b111100000000;
20'b01101001110101111111: color_data = 12'b111100000000;
20'b01101001110110000000: color_data = 12'b111100000000;
20'b01101001110110000001: color_data = 12'b111100000000;
20'b01101001110110000010: color_data = 12'b111100000000;
20'b01101001110110000011: color_data = 12'b111100000000;
20'b01101001110110000100: color_data = 12'b111100000000;
20'b01101001110110000101: color_data = 12'b111100000000;
20'b01101001110110000110: color_data = 12'b111100000000;
20'b01101001110110000111: color_data = 12'b111100000000;
20'b01101001110110001000: color_data = 12'b111100000000;
20'b01101001110110001001: color_data = 12'b111100000000;
20'b01101001110110001101: color_data = 12'b111100000000;
20'b01101001110110001110: color_data = 12'b111100000000;
20'b01101001110110001111: color_data = 12'b111100000000;
20'b01101001110110010000: color_data = 12'b111100000000;
20'b01101001110110010001: color_data = 12'b111100000000;
20'b01101001110110010010: color_data = 12'b111100000000;
20'b01101001110110010011: color_data = 12'b111100000000;
20'b01101001110110010100: color_data = 12'b111100000000;
20'b01101001110110010101: color_data = 12'b111100000000;
20'b01101001110110010110: color_data = 12'b111100000000;
20'b01101001110110010111: color_data = 12'b111100000000;
20'b01101001110110011000: color_data = 12'b111100000000;
20'b01101001110110011001: color_data = 12'b111100000000;
20'b01101001110110011010: color_data = 12'b111100000000;
20'b01101001110110011011: color_data = 12'b111100000000;
20'b01101001110110011100: color_data = 12'b111100000000;
20'b01101001110110011101: color_data = 12'b111100000000;
20'b01101001110110011110: color_data = 12'b111100000000;
20'b01101010000011111010: color_data = 12'b111101110000;
20'b01101010000011111011: color_data = 12'b111101110000;
20'b01101010000011111100: color_data = 12'b111101110000;
20'b01101010000011111101: color_data = 12'b111101110000;
20'b01101010000011111110: color_data = 12'b111101110000;
20'b01101010000011111111: color_data = 12'b111101110000;
20'b01101010000100000000: color_data = 12'b111101110000;
20'b01101010000100000001: color_data = 12'b111101110000;
20'b01101010000100000010: color_data = 12'b111101110000;
20'b01101010000100000011: color_data = 12'b111101110000;
20'b01101010000100000100: color_data = 12'b111101110000;
20'b01101010000100000101: color_data = 12'b111101110000;
20'b01101010000100000110: color_data = 12'b111101110000;
20'b01101010000100000111: color_data = 12'b111101110000;
20'b01101010000100001000: color_data = 12'b111101110000;
20'b01101010000100001001: color_data = 12'b111101110000;
20'b01101010000100001010: color_data = 12'b111101110000;
20'b01101010000100001011: color_data = 12'b111101110000;
20'b01101010000100001111: color_data = 12'b111101110000;
20'b01101010000100010000: color_data = 12'b111101110000;
20'b01101010000100010001: color_data = 12'b111101110000;
20'b01101010000100010010: color_data = 12'b111101110000;
20'b01101010000100010011: color_data = 12'b111101110000;
20'b01101010000100010100: color_data = 12'b111101110000;
20'b01101010000100010101: color_data = 12'b111101110000;
20'b01101010000100010110: color_data = 12'b111101110000;
20'b01101010000100010111: color_data = 12'b111101110000;
20'b01101010000100011000: color_data = 12'b111101110000;
20'b01101010000100011001: color_data = 12'b111101110000;
20'b01101010000100011010: color_data = 12'b111101110000;
20'b01101010000100011011: color_data = 12'b111101110000;
20'b01101010000100011100: color_data = 12'b111101110000;
20'b01101010000100011101: color_data = 12'b111101110000;
20'b01101010000100011110: color_data = 12'b111101110000;
20'b01101010000100011111: color_data = 12'b111101110000;
20'b01101010000100100000: color_data = 12'b111101110000;
20'b01101010000100100100: color_data = 12'b111101110000;
20'b01101010000100100101: color_data = 12'b111101110000;
20'b01101010000100100110: color_data = 12'b111101110000;
20'b01101010000100100111: color_data = 12'b111101110000;
20'b01101010000100101000: color_data = 12'b111101110000;
20'b01101010000100101001: color_data = 12'b111101110000;
20'b01101010000100101010: color_data = 12'b111101110000;
20'b01101010000100101011: color_data = 12'b111101110000;
20'b01101010000100101100: color_data = 12'b111101110000;
20'b01101010000100101101: color_data = 12'b111101110000;
20'b01101010000100101110: color_data = 12'b111101110000;
20'b01101010000100101111: color_data = 12'b111101110000;
20'b01101010000100110000: color_data = 12'b111101110000;
20'b01101010000100110001: color_data = 12'b111101110000;
20'b01101010000100110010: color_data = 12'b111101110000;
20'b01101010000100110011: color_data = 12'b111101110000;
20'b01101010000100110100: color_data = 12'b111101110000;
20'b01101010000100110101: color_data = 12'b111101110000;
20'b01101010000100111001: color_data = 12'b111101110000;
20'b01101010000100111010: color_data = 12'b111101110000;
20'b01101010000100111011: color_data = 12'b111101110000;
20'b01101010000100111100: color_data = 12'b111101110000;
20'b01101010000100111101: color_data = 12'b111101110000;
20'b01101010000100111110: color_data = 12'b111101110000;
20'b01101010000100111111: color_data = 12'b111101110000;
20'b01101010000101000000: color_data = 12'b111101110000;
20'b01101010000101000001: color_data = 12'b111101110000;
20'b01101010000101000010: color_data = 12'b111101110000;
20'b01101010000101000011: color_data = 12'b111101110000;
20'b01101010000101000100: color_data = 12'b111101110000;
20'b01101010000101000101: color_data = 12'b111101110000;
20'b01101010000101000110: color_data = 12'b111101110000;
20'b01101010000101000111: color_data = 12'b111101110000;
20'b01101010000101001000: color_data = 12'b111101110000;
20'b01101010000101001001: color_data = 12'b111101110000;
20'b01101010000101001010: color_data = 12'b111101110000;
20'b01101010000101001110: color_data = 12'b000011110000;
20'b01101010000101001111: color_data = 12'b000011110000;
20'b01101010000101010000: color_data = 12'b000011110000;
20'b01101010000101010001: color_data = 12'b000011110000;
20'b01101010000101010010: color_data = 12'b000011110000;
20'b01101010000101010011: color_data = 12'b000011110000;
20'b01101010000101010100: color_data = 12'b000011110000;
20'b01101010000101010101: color_data = 12'b000011110000;
20'b01101010000101010110: color_data = 12'b000011110000;
20'b01101010000101010111: color_data = 12'b000011110000;
20'b01101010000101011000: color_data = 12'b000011110000;
20'b01101010000101011001: color_data = 12'b000011110000;
20'b01101010000101011010: color_data = 12'b000011110000;
20'b01101010000101011011: color_data = 12'b000011110000;
20'b01101010000101011100: color_data = 12'b000011110000;
20'b01101010000101011101: color_data = 12'b000011110000;
20'b01101010000101011110: color_data = 12'b000011110000;
20'b01101010000101011111: color_data = 12'b000011110000;
20'b01101010000101100011: color_data = 12'b111100001111;
20'b01101010000101100100: color_data = 12'b111100001111;
20'b01101010000101100101: color_data = 12'b111100001111;
20'b01101010000101100110: color_data = 12'b111100001111;
20'b01101010000101100111: color_data = 12'b111100001111;
20'b01101010000101101000: color_data = 12'b111100001111;
20'b01101010000101101001: color_data = 12'b111100001111;
20'b01101010000101101010: color_data = 12'b111100001111;
20'b01101010000101101011: color_data = 12'b111100001111;
20'b01101010000101101100: color_data = 12'b111100001111;
20'b01101010000101101101: color_data = 12'b111100001111;
20'b01101010000101101110: color_data = 12'b111100001111;
20'b01101010000101101111: color_data = 12'b111100001111;
20'b01101010000101110000: color_data = 12'b111100001111;
20'b01101010000101110001: color_data = 12'b111100001111;
20'b01101010000101110010: color_data = 12'b111100001111;
20'b01101010000101110011: color_data = 12'b111100001111;
20'b01101010000101110100: color_data = 12'b111100001111;
20'b01101010000101111000: color_data = 12'b111100000000;
20'b01101010000101111001: color_data = 12'b111100000000;
20'b01101010000101111010: color_data = 12'b111100000000;
20'b01101010000101111011: color_data = 12'b111100000000;
20'b01101010000101111100: color_data = 12'b111100000000;
20'b01101010000101111101: color_data = 12'b111100000000;
20'b01101010000101111110: color_data = 12'b111100000000;
20'b01101010000101111111: color_data = 12'b111100000000;
20'b01101010000110000000: color_data = 12'b111100000000;
20'b01101010000110000001: color_data = 12'b111100000000;
20'b01101010000110000010: color_data = 12'b111100000000;
20'b01101010000110000011: color_data = 12'b111100000000;
20'b01101010000110000100: color_data = 12'b111100000000;
20'b01101010000110000101: color_data = 12'b111100000000;
20'b01101010000110000110: color_data = 12'b111100000000;
20'b01101010000110000111: color_data = 12'b111100000000;
20'b01101010000110001000: color_data = 12'b111100000000;
20'b01101010000110001001: color_data = 12'b111100000000;
20'b01101010000110001101: color_data = 12'b111100000000;
20'b01101010000110001110: color_data = 12'b111100000000;
20'b01101010000110001111: color_data = 12'b111100000000;
20'b01101010000110010000: color_data = 12'b111100000000;
20'b01101010000110010001: color_data = 12'b111100000000;
20'b01101010000110010010: color_data = 12'b111100000000;
20'b01101010000110010011: color_data = 12'b111100000000;
20'b01101010000110010100: color_data = 12'b111100000000;
20'b01101010000110010101: color_data = 12'b111100000000;
20'b01101010000110010110: color_data = 12'b111100000000;
20'b01101010000110010111: color_data = 12'b111100000000;
20'b01101010000110011000: color_data = 12'b111100000000;
20'b01101010000110011001: color_data = 12'b111100000000;
20'b01101010000110011010: color_data = 12'b111100000000;
20'b01101010000110011011: color_data = 12'b111100000000;
20'b01101010000110011100: color_data = 12'b111100000000;
20'b01101010000110011101: color_data = 12'b111100000000;
20'b01101010000110011110: color_data = 12'b111100000000;
20'b01101010010011111010: color_data = 12'b111101110000;
20'b01101010010011111011: color_data = 12'b111101110000;
20'b01101010010011111100: color_data = 12'b111101110000;
20'b01101010010011111101: color_data = 12'b111101110000;
20'b01101010010011111110: color_data = 12'b111101110000;
20'b01101010010011111111: color_data = 12'b111101110000;
20'b01101010010100000000: color_data = 12'b111101110000;
20'b01101010010100000001: color_data = 12'b111101110000;
20'b01101010010100000010: color_data = 12'b111101110000;
20'b01101010010100000011: color_data = 12'b111101110000;
20'b01101010010100000100: color_data = 12'b111101110000;
20'b01101010010100000101: color_data = 12'b111101110000;
20'b01101010010100000110: color_data = 12'b111101110000;
20'b01101010010100000111: color_data = 12'b111101110000;
20'b01101010010100001000: color_data = 12'b111101110000;
20'b01101010010100001001: color_data = 12'b111101110000;
20'b01101010010100001010: color_data = 12'b111101110000;
20'b01101010010100001011: color_data = 12'b111101110000;
20'b01101010010100001111: color_data = 12'b111101110000;
20'b01101010010100010000: color_data = 12'b111101110000;
20'b01101010010100010001: color_data = 12'b111101110000;
20'b01101010010100010010: color_data = 12'b111101110000;
20'b01101010010100010011: color_data = 12'b111101110000;
20'b01101010010100010100: color_data = 12'b111101110000;
20'b01101010010100010101: color_data = 12'b111101110000;
20'b01101010010100010110: color_data = 12'b111101110000;
20'b01101010010100010111: color_data = 12'b111101110000;
20'b01101010010100011000: color_data = 12'b111101110000;
20'b01101010010100011001: color_data = 12'b111101110000;
20'b01101010010100011010: color_data = 12'b111101110000;
20'b01101010010100011011: color_data = 12'b111101110000;
20'b01101010010100011100: color_data = 12'b111101110000;
20'b01101010010100011101: color_data = 12'b111101110000;
20'b01101010010100011110: color_data = 12'b111101110000;
20'b01101010010100011111: color_data = 12'b111101110000;
20'b01101010010100100000: color_data = 12'b111101110000;
20'b01101010010100100100: color_data = 12'b111101110000;
20'b01101010010100100101: color_data = 12'b111101110000;
20'b01101010010100100110: color_data = 12'b111101110000;
20'b01101010010100100111: color_data = 12'b111101110000;
20'b01101010010100101000: color_data = 12'b111101110000;
20'b01101010010100101001: color_data = 12'b111101110000;
20'b01101010010100101010: color_data = 12'b111101110000;
20'b01101010010100101011: color_data = 12'b111101110000;
20'b01101010010100101100: color_data = 12'b111101110000;
20'b01101010010100101101: color_data = 12'b111101110000;
20'b01101010010100101110: color_data = 12'b111101110000;
20'b01101010010100101111: color_data = 12'b111101110000;
20'b01101010010100110000: color_data = 12'b111101110000;
20'b01101010010100110001: color_data = 12'b111101110000;
20'b01101010010100110010: color_data = 12'b111101110000;
20'b01101010010100110011: color_data = 12'b111101110000;
20'b01101010010100110100: color_data = 12'b111101110000;
20'b01101010010100110101: color_data = 12'b111101110000;
20'b01101010010100111001: color_data = 12'b111101110000;
20'b01101010010100111010: color_data = 12'b111101110000;
20'b01101010010100111011: color_data = 12'b111101110000;
20'b01101010010100111100: color_data = 12'b111101110000;
20'b01101010010100111101: color_data = 12'b111101110000;
20'b01101010010100111110: color_data = 12'b111101110000;
20'b01101010010100111111: color_data = 12'b111101110000;
20'b01101010010101000000: color_data = 12'b111101110000;
20'b01101010010101000001: color_data = 12'b111101110000;
20'b01101010010101000010: color_data = 12'b111101110000;
20'b01101010010101000011: color_data = 12'b111101110000;
20'b01101010010101000100: color_data = 12'b111101110000;
20'b01101010010101000101: color_data = 12'b111101110000;
20'b01101010010101000110: color_data = 12'b111101110000;
20'b01101010010101000111: color_data = 12'b111101110000;
20'b01101010010101001000: color_data = 12'b111101110000;
20'b01101010010101001001: color_data = 12'b111101110000;
20'b01101010010101001010: color_data = 12'b111101110000;
20'b01101010010101001110: color_data = 12'b000011110000;
20'b01101010010101001111: color_data = 12'b000011110000;
20'b01101010010101010000: color_data = 12'b000011110000;
20'b01101010010101010001: color_data = 12'b000011110000;
20'b01101010010101010010: color_data = 12'b000011110000;
20'b01101010010101010011: color_data = 12'b000011110000;
20'b01101010010101010100: color_data = 12'b000011110000;
20'b01101010010101010101: color_data = 12'b000011110000;
20'b01101010010101010110: color_data = 12'b000011110000;
20'b01101010010101010111: color_data = 12'b000011110000;
20'b01101010010101011000: color_data = 12'b000011110000;
20'b01101010010101011001: color_data = 12'b000011110000;
20'b01101010010101011010: color_data = 12'b000011110000;
20'b01101010010101011011: color_data = 12'b000011110000;
20'b01101010010101011100: color_data = 12'b000011110000;
20'b01101010010101011101: color_data = 12'b000011110000;
20'b01101010010101011110: color_data = 12'b000011110000;
20'b01101010010101011111: color_data = 12'b000011110000;
20'b01101010010101100011: color_data = 12'b111100001111;
20'b01101010010101100100: color_data = 12'b111100001111;
20'b01101010010101100101: color_data = 12'b111100001111;
20'b01101010010101100110: color_data = 12'b111100001111;
20'b01101010010101100111: color_data = 12'b111100001111;
20'b01101010010101101000: color_data = 12'b111100001111;
20'b01101010010101101001: color_data = 12'b111100001111;
20'b01101010010101101010: color_data = 12'b111100001111;
20'b01101010010101101011: color_data = 12'b111100001111;
20'b01101010010101101100: color_data = 12'b111100001111;
20'b01101010010101101101: color_data = 12'b111100001111;
20'b01101010010101101110: color_data = 12'b111100001111;
20'b01101010010101101111: color_data = 12'b111100001111;
20'b01101010010101110000: color_data = 12'b111100001111;
20'b01101010010101110001: color_data = 12'b111100001111;
20'b01101010010101110010: color_data = 12'b111100001111;
20'b01101010010101110011: color_data = 12'b111100001111;
20'b01101010010101110100: color_data = 12'b111100001111;
20'b01101010010101111000: color_data = 12'b111100000000;
20'b01101010010101111001: color_data = 12'b111100000000;
20'b01101010010101111010: color_data = 12'b111100000000;
20'b01101010010101111011: color_data = 12'b111100000000;
20'b01101010010101111100: color_data = 12'b111100000000;
20'b01101010010101111101: color_data = 12'b111100000000;
20'b01101010010101111110: color_data = 12'b111100000000;
20'b01101010010101111111: color_data = 12'b111100000000;
20'b01101010010110000000: color_data = 12'b111100000000;
20'b01101010010110000001: color_data = 12'b111100000000;
20'b01101010010110000010: color_data = 12'b111100000000;
20'b01101010010110000011: color_data = 12'b111100000000;
20'b01101010010110000100: color_data = 12'b111100000000;
20'b01101010010110000101: color_data = 12'b111100000000;
20'b01101010010110000110: color_data = 12'b111100000000;
20'b01101010010110000111: color_data = 12'b111100000000;
20'b01101010010110001000: color_data = 12'b111100000000;
20'b01101010010110001001: color_data = 12'b111100000000;
20'b01101010010110001101: color_data = 12'b111100000000;
20'b01101010010110001110: color_data = 12'b111100000000;
20'b01101010010110001111: color_data = 12'b111100000000;
20'b01101010010110010000: color_data = 12'b111100000000;
20'b01101010010110010001: color_data = 12'b111100000000;
20'b01101010010110010010: color_data = 12'b111100000000;
20'b01101010010110010011: color_data = 12'b111100000000;
20'b01101010010110010100: color_data = 12'b111100000000;
20'b01101010010110010101: color_data = 12'b111100000000;
20'b01101010010110010110: color_data = 12'b111100000000;
20'b01101010010110010111: color_data = 12'b111100000000;
20'b01101010010110011000: color_data = 12'b111100000000;
20'b01101010010110011001: color_data = 12'b111100000000;
20'b01101010010110011010: color_data = 12'b111100000000;
20'b01101010010110011011: color_data = 12'b111100000000;
20'b01101010010110011100: color_data = 12'b111100000000;
20'b01101010010110011101: color_data = 12'b111100000000;
20'b01101010010110011110: color_data = 12'b111100000000;
20'b01101010100011111010: color_data = 12'b111101110000;
20'b01101010100011111011: color_data = 12'b111101110000;
20'b01101010100011111100: color_data = 12'b111101110000;
20'b01101010100011111101: color_data = 12'b111101110000;
20'b01101010100011111110: color_data = 12'b111101110000;
20'b01101010100011111111: color_data = 12'b111101110000;
20'b01101010100100000000: color_data = 12'b111101110000;
20'b01101010100100000001: color_data = 12'b111101110000;
20'b01101010100100000010: color_data = 12'b111101110000;
20'b01101010100100000011: color_data = 12'b111101110000;
20'b01101010100100000100: color_data = 12'b111101110000;
20'b01101010100100000101: color_data = 12'b111101110000;
20'b01101010100100000110: color_data = 12'b111101110000;
20'b01101010100100000111: color_data = 12'b111101110000;
20'b01101010100100001000: color_data = 12'b111101110000;
20'b01101010100100001001: color_data = 12'b111101110000;
20'b01101010100100001010: color_data = 12'b111101110000;
20'b01101010100100001011: color_data = 12'b111101110000;
20'b01101010100100001111: color_data = 12'b111101110000;
20'b01101010100100010000: color_data = 12'b111101110000;
20'b01101010100100010001: color_data = 12'b111101110000;
20'b01101010100100010010: color_data = 12'b111101110000;
20'b01101010100100010011: color_data = 12'b111101110000;
20'b01101010100100010100: color_data = 12'b111101110000;
20'b01101010100100010101: color_data = 12'b111101110000;
20'b01101010100100010110: color_data = 12'b111101110000;
20'b01101010100100010111: color_data = 12'b111101110000;
20'b01101010100100011000: color_data = 12'b111101110000;
20'b01101010100100011001: color_data = 12'b111101110000;
20'b01101010100100011010: color_data = 12'b111101110000;
20'b01101010100100011011: color_data = 12'b111101110000;
20'b01101010100100011100: color_data = 12'b111101110000;
20'b01101010100100011101: color_data = 12'b111101110000;
20'b01101010100100011110: color_data = 12'b111101110000;
20'b01101010100100011111: color_data = 12'b111101110000;
20'b01101010100100100000: color_data = 12'b111101110000;
20'b01101010100100100100: color_data = 12'b111101110000;
20'b01101010100100100101: color_data = 12'b111101110000;
20'b01101010100100100110: color_data = 12'b111101110000;
20'b01101010100100100111: color_data = 12'b111101110000;
20'b01101010100100101000: color_data = 12'b111101110000;
20'b01101010100100101001: color_data = 12'b111101110000;
20'b01101010100100101010: color_data = 12'b111101110000;
20'b01101010100100101011: color_data = 12'b111101110000;
20'b01101010100100101100: color_data = 12'b111101110000;
20'b01101010100100101101: color_data = 12'b111101110000;
20'b01101010100100101110: color_data = 12'b111101110000;
20'b01101010100100101111: color_data = 12'b111101110000;
20'b01101010100100110000: color_data = 12'b111101110000;
20'b01101010100100110001: color_data = 12'b111101110000;
20'b01101010100100110010: color_data = 12'b111101110000;
20'b01101010100100110011: color_data = 12'b111101110000;
20'b01101010100100110100: color_data = 12'b111101110000;
20'b01101010100100110101: color_data = 12'b111101110000;
20'b01101010100100111001: color_data = 12'b111101110000;
20'b01101010100100111010: color_data = 12'b111101110000;
20'b01101010100100111011: color_data = 12'b111101110000;
20'b01101010100100111100: color_data = 12'b111101110000;
20'b01101010100100111101: color_data = 12'b111101110000;
20'b01101010100100111110: color_data = 12'b111101110000;
20'b01101010100100111111: color_data = 12'b111101110000;
20'b01101010100101000000: color_data = 12'b111101110000;
20'b01101010100101000001: color_data = 12'b111101110000;
20'b01101010100101000010: color_data = 12'b111101110000;
20'b01101010100101000011: color_data = 12'b111101110000;
20'b01101010100101000100: color_data = 12'b111101110000;
20'b01101010100101000101: color_data = 12'b111101110000;
20'b01101010100101000110: color_data = 12'b111101110000;
20'b01101010100101000111: color_data = 12'b111101110000;
20'b01101010100101001000: color_data = 12'b111101110000;
20'b01101010100101001001: color_data = 12'b111101110000;
20'b01101010100101001010: color_data = 12'b111101110000;
20'b01101010100101001110: color_data = 12'b000011110000;
20'b01101010100101001111: color_data = 12'b000011110000;
20'b01101010100101010000: color_data = 12'b000011110000;
20'b01101010100101010001: color_data = 12'b000011110000;
20'b01101010100101010010: color_data = 12'b000011110000;
20'b01101010100101010011: color_data = 12'b000011110000;
20'b01101010100101010100: color_data = 12'b000011110000;
20'b01101010100101010101: color_data = 12'b000011110000;
20'b01101010100101010110: color_data = 12'b000011110000;
20'b01101010100101010111: color_data = 12'b000011110000;
20'b01101010100101011000: color_data = 12'b000011110000;
20'b01101010100101011001: color_data = 12'b000011110000;
20'b01101010100101011010: color_data = 12'b000011110000;
20'b01101010100101011011: color_data = 12'b000011110000;
20'b01101010100101011100: color_data = 12'b000011110000;
20'b01101010100101011101: color_data = 12'b000011110000;
20'b01101010100101011110: color_data = 12'b000011110000;
20'b01101010100101011111: color_data = 12'b000011110000;
20'b01101010100101100011: color_data = 12'b111100001111;
20'b01101010100101100100: color_data = 12'b111100001111;
20'b01101010100101100101: color_data = 12'b111100001111;
20'b01101010100101100110: color_data = 12'b111100001111;
20'b01101010100101100111: color_data = 12'b111100001111;
20'b01101010100101101000: color_data = 12'b111100001111;
20'b01101010100101101001: color_data = 12'b111100001111;
20'b01101010100101101010: color_data = 12'b111100001111;
20'b01101010100101101011: color_data = 12'b111100001111;
20'b01101010100101101100: color_data = 12'b111100001111;
20'b01101010100101101101: color_data = 12'b111100001111;
20'b01101010100101101110: color_data = 12'b111100001111;
20'b01101010100101101111: color_data = 12'b111100001111;
20'b01101010100101110000: color_data = 12'b111100001111;
20'b01101010100101110001: color_data = 12'b111100001111;
20'b01101010100101110010: color_data = 12'b111100001111;
20'b01101010100101110011: color_data = 12'b111100001111;
20'b01101010100101110100: color_data = 12'b111100001111;
20'b01101010100101111000: color_data = 12'b111100000000;
20'b01101010100101111001: color_data = 12'b111100000000;
20'b01101010100101111010: color_data = 12'b111100000000;
20'b01101010100101111011: color_data = 12'b111100000000;
20'b01101010100101111100: color_data = 12'b111100000000;
20'b01101010100101111101: color_data = 12'b111100000000;
20'b01101010100101111110: color_data = 12'b111100000000;
20'b01101010100101111111: color_data = 12'b111100000000;
20'b01101010100110000000: color_data = 12'b111100000000;
20'b01101010100110000001: color_data = 12'b111100000000;
20'b01101010100110000010: color_data = 12'b111100000000;
20'b01101010100110000011: color_data = 12'b111100000000;
20'b01101010100110000100: color_data = 12'b111100000000;
20'b01101010100110000101: color_data = 12'b111100000000;
20'b01101010100110000110: color_data = 12'b111100000000;
20'b01101010100110000111: color_data = 12'b111100000000;
20'b01101010100110001000: color_data = 12'b111100000000;
20'b01101010100110001001: color_data = 12'b111100000000;
20'b01101010100110001101: color_data = 12'b111100000000;
20'b01101010100110001110: color_data = 12'b111100000000;
20'b01101010100110001111: color_data = 12'b111100000000;
20'b01101010100110010000: color_data = 12'b111100000000;
20'b01101010100110010001: color_data = 12'b111100000000;
20'b01101010100110010010: color_data = 12'b111100000000;
20'b01101010100110010011: color_data = 12'b111100000000;
20'b01101010100110010100: color_data = 12'b111100000000;
20'b01101010100110010101: color_data = 12'b111100000000;
20'b01101010100110010110: color_data = 12'b111100000000;
20'b01101010100110010111: color_data = 12'b111100000000;
20'b01101010100110011000: color_data = 12'b111100000000;
20'b01101010100110011001: color_data = 12'b111100000000;
20'b01101010100110011010: color_data = 12'b111100000000;
20'b01101010100110011011: color_data = 12'b111100000000;
20'b01101010100110011100: color_data = 12'b111100000000;
20'b01101010100110011101: color_data = 12'b111100000000;
20'b01101010100110011110: color_data = 12'b111100000000;
20'b01101010110011111010: color_data = 12'b111101110000;
20'b01101010110011111011: color_data = 12'b111101110000;
20'b01101010110011111100: color_data = 12'b111101110000;
20'b01101010110011111101: color_data = 12'b111101110000;
20'b01101010110011111110: color_data = 12'b111101110000;
20'b01101010110011111111: color_data = 12'b111101110000;
20'b01101010110100000000: color_data = 12'b111101110000;
20'b01101010110100000001: color_data = 12'b111101110000;
20'b01101010110100000010: color_data = 12'b111101110000;
20'b01101010110100000011: color_data = 12'b111101110000;
20'b01101010110100000100: color_data = 12'b111101110000;
20'b01101010110100000101: color_data = 12'b111101110000;
20'b01101010110100000110: color_data = 12'b111101110000;
20'b01101010110100000111: color_data = 12'b111101110000;
20'b01101010110100001000: color_data = 12'b111101110000;
20'b01101010110100001001: color_data = 12'b111101110000;
20'b01101010110100001010: color_data = 12'b111101110000;
20'b01101010110100001011: color_data = 12'b111101110000;
20'b01101010110100001111: color_data = 12'b111101110000;
20'b01101010110100010000: color_data = 12'b111101110000;
20'b01101010110100010001: color_data = 12'b111101110000;
20'b01101010110100010010: color_data = 12'b111101110000;
20'b01101010110100010011: color_data = 12'b111101110000;
20'b01101010110100010100: color_data = 12'b111101110000;
20'b01101010110100010101: color_data = 12'b111101110000;
20'b01101010110100010110: color_data = 12'b111101110000;
20'b01101010110100010111: color_data = 12'b111101110000;
20'b01101010110100011000: color_data = 12'b111101110000;
20'b01101010110100011001: color_data = 12'b111101110000;
20'b01101010110100011010: color_data = 12'b111101110000;
20'b01101010110100011011: color_data = 12'b111101110000;
20'b01101010110100011100: color_data = 12'b111101110000;
20'b01101010110100011101: color_data = 12'b111101110000;
20'b01101010110100011110: color_data = 12'b111101110000;
20'b01101010110100011111: color_data = 12'b111101110000;
20'b01101010110100100000: color_data = 12'b111101110000;
20'b01101010110100100100: color_data = 12'b111101110000;
20'b01101010110100100101: color_data = 12'b111101110000;
20'b01101010110100100110: color_data = 12'b111101110000;
20'b01101010110100100111: color_data = 12'b111101110000;
20'b01101010110100101000: color_data = 12'b111101110000;
20'b01101010110100101001: color_data = 12'b111101110000;
20'b01101010110100101010: color_data = 12'b111101110000;
20'b01101010110100101011: color_data = 12'b111101110000;
20'b01101010110100101100: color_data = 12'b111101110000;
20'b01101010110100101101: color_data = 12'b111101110000;
20'b01101010110100101110: color_data = 12'b111101110000;
20'b01101010110100101111: color_data = 12'b111101110000;
20'b01101010110100110000: color_data = 12'b111101110000;
20'b01101010110100110001: color_data = 12'b111101110000;
20'b01101010110100110010: color_data = 12'b111101110000;
20'b01101010110100110011: color_data = 12'b111101110000;
20'b01101010110100110100: color_data = 12'b111101110000;
20'b01101010110100110101: color_data = 12'b111101110000;
20'b01101010110100111001: color_data = 12'b111101110000;
20'b01101010110100111010: color_data = 12'b111101110000;
20'b01101010110100111011: color_data = 12'b111101110000;
20'b01101010110100111100: color_data = 12'b111101110000;
20'b01101010110100111101: color_data = 12'b111101110000;
20'b01101010110100111110: color_data = 12'b111101110000;
20'b01101010110100111111: color_data = 12'b111101110000;
20'b01101010110101000000: color_data = 12'b111101110000;
20'b01101010110101000001: color_data = 12'b111101110000;
20'b01101010110101000010: color_data = 12'b111101110000;
20'b01101010110101000011: color_data = 12'b111101110000;
20'b01101010110101000100: color_data = 12'b111101110000;
20'b01101010110101000101: color_data = 12'b111101110000;
20'b01101010110101000110: color_data = 12'b111101110000;
20'b01101010110101000111: color_data = 12'b111101110000;
20'b01101010110101001000: color_data = 12'b111101110000;
20'b01101010110101001001: color_data = 12'b111101110000;
20'b01101010110101001010: color_data = 12'b111101110000;
20'b01101010110101001110: color_data = 12'b000011110000;
20'b01101010110101001111: color_data = 12'b000011110000;
20'b01101010110101010000: color_data = 12'b000011110000;
20'b01101010110101010001: color_data = 12'b000011110000;
20'b01101010110101010010: color_data = 12'b000011110000;
20'b01101010110101010011: color_data = 12'b000011110000;
20'b01101010110101010100: color_data = 12'b000011110000;
20'b01101010110101010101: color_data = 12'b000011110000;
20'b01101010110101010110: color_data = 12'b000011110000;
20'b01101010110101010111: color_data = 12'b000011110000;
20'b01101010110101011000: color_data = 12'b000011110000;
20'b01101010110101011001: color_data = 12'b000011110000;
20'b01101010110101011010: color_data = 12'b000011110000;
20'b01101010110101011011: color_data = 12'b000011110000;
20'b01101010110101011100: color_data = 12'b000011110000;
20'b01101010110101011101: color_data = 12'b000011110000;
20'b01101010110101011110: color_data = 12'b000011110000;
20'b01101010110101011111: color_data = 12'b000011110000;
20'b01101010110101100011: color_data = 12'b111100001111;
20'b01101010110101100100: color_data = 12'b111100001111;
20'b01101010110101100101: color_data = 12'b111100001111;
20'b01101010110101100110: color_data = 12'b111100001111;
20'b01101010110101100111: color_data = 12'b111100001111;
20'b01101010110101101000: color_data = 12'b111100001111;
20'b01101010110101101001: color_data = 12'b111100001111;
20'b01101010110101101010: color_data = 12'b111100001111;
20'b01101010110101101011: color_data = 12'b111100001111;
20'b01101010110101101100: color_data = 12'b111100001111;
20'b01101010110101101101: color_data = 12'b111100001111;
20'b01101010110101101110: color_data = 12'b111100001111;
20'b01101010110101101111: color_data = 12'b111100001111;
20'b01101010110101110000: color_data = 12'b111100001111;
20'b01101010110101110001: color_data = 12'b111100001111;
20'b01101010110101110010: color_data = 12'b111100001111;
20'b01101010110101110011: color_data = 12'b111100001111;
20'b01101010110101110100: color_data = 12'b111100001111;
20'b01101010110101111000: color_data = 12'b111100000000;
20'b01101010110101111001: color_data = 12'b111100000000;
20'b01101010110101111010: color_data = 12'b111100000000;
20'b01101010110101111011: color_data = 12'b111100000000;
20'b01101010110101111100: color_data = 12'b111100000000;
20'b01101010110101111101: color_data = 12'b111100000000;
20'b01101010110101111110: color_data = 12'b111100000000;
20'b01101010110101111111: color_data = 12'b111100000000;
20'b01101010110110000000: color_data = 12'b111100000000;
20'b01101010110110000001: color_data = 12'b111100000000;
20'b01101010110110000010: color_data = 12'b111100000000;
20'b01101010110110000011: color_data = 12'b111100000000;
20'b01101010110110000100: color_data = 12'b111100000000;
20'b01101010110110000101: color_data = 12'b111100000000;
20'b01101010110110000110: color_data = 12'b111100000000;
20'b01101010110110000111: color_data = 12'b111100000000;
20'b01101010110110001000: color_data = 12'b111100000000;
20'b01101010110110001001: color_data = 12'b111100000000;
20'b01101010110110001101: color_data = 12'b111100000000;
20'b01101010110110001110: color_data = 12'b111100000000;
20'b01101010110110001111: color_data = 12'b111100000000;
20'b01101010110110010000: color_data = 12'b111100000000;
20'b01101010110110010001: color_data = 12'b111100000000;
20'b01101010110110010010: color_data = 12'b111100000000;
20'b01101010110110010011: color_data = 12'b111100000000;
20'b01101010110110010100: color_data = 12'b111100000000;
20'b01101010110110010101: color_data = 12'b111100000000;
20'b01101010110110010110: color_data = 12'b111100000000;
20'b01101010110110010111: color_data = 12'b111100000000;
20'b01101010110110011000: color_data = 12'b111100000000;
20'b01101010110110011001: color_data = 12'b111100000000;
20'b01101010110110011010: color_data = 12'b111100000000;
20'b01101010110110011011: color_data = 12'b111100000000;
20'b01101010110110011100: color_data = 12'b111100000000;
20'b01101010110110011101: color_data = 12'b111100000000;
20'b01101010110110011110: color_data = 12'b111100000000;
20'b01101011000011111010: color_data = 12'b111101110000;
20'b01101011000011111011: color_data = 12'b111101110000;
20'b01101011000011111100: color_data = 12'b111101110000;
20'b01101011000011111101: color_data = 12'b111101110000;
20'b01101011000011111110: color_data = 12'b111101110000;
20'b01101011000011111111: color_data = 12'b111101110000;
20'b01101011000100000000: color_data = 12'b111101110000;
20'b01101011000100000001: color_data = 12'b111101110000;
20'b01101011000100000010: color_data = 12'b111101110000;
20'b01101011000100000011: color_data = 12'b111101110000;
20'b01101011000100000100: color_data = 12'b111101110000;
20'b01101011000100000101: color_data = 12'b111101110000;
20'b01101011000100000110: color_data = 12'b111101110000;
20'b01101011000100000111: color_data = 12'b111101110000;
20'b01101011000100001000: color_data = 12'b111101110000;
20'b01101011000100001001: color_data = 12'b111101110000;
20'b01101011000100001010: color_data = 12'b111101110000;
20'b01101011000100001011: color_data = 12'b111101110000;
20'b01101011000100001111: color_data = 12'b111101110000;
20'b01101011000100010000: color_data = 12'b111101110000;
20'b01101011000100010001: color_data = 12'b111101110000;
20'b01101011000100010010: color_data = 12'b111101110000;
20'b01101011000100010011: color_data = 12'b111101110000;
20'b01101011000100010100: color_data = 12'b111101110000;
20'b01101011000100010101: color_data = 12'b111101110000;
20'b01101011000100010110: color_data = 12'b111101110000;
20'b01101011000100010111: color_data = 12'b111101110000;
20'b01101011000100011000: color_data = 12'b111101110000;
20'b01101011000100011001: color_data = 12'b111101110000;
20'b01101011000100011010: color_data = 12'b111101110000;
20'b01101011000100011011: color_data = 12'b111101110000;
20'b01101011000100011100: color_data = 12'b111101110000;
20'b01101011000100011101: color_data = 12'b111101110000;
20'b01101011000100011110: color_data = 12'b111101110000;
20'b01101011000100011111: color_data = 12'b111101110000;
20'b01101011000100100000: color_data = 12'b111101110000;
20'b01101011000100100100: color_data = 12'b111101110000;
20'b01101011000100100101: color_data = 12'b111101110000;
20'b01101011000100100110: color_data = 12'b111101110000;
20'b01101011000100100111: color_data = 12'b111101110000;
20'b01101011000100101000: color_data = 12'b111101110000;
20'b01101011000100101001: color_data = 12'b111101110000;
20'b01101011000100101010: color_data = 12'b111101110000;
20'b01101011000100101011: color_data = 12'b111101110000;
20'b01101011000100101100: color_data = 12'b111101110000;
20'b01101011000100101101: color_data = 12'b111101110000;
20'b01101011000100101110: color_data = 12'b111101110000;
20'b01101011000100101111: color_data = 12'b111101110000;
20'b01101011000100110000: color_data = 12'b111101110000;
20'b01101011000100110001: color_data = 12'b111101110000;
20'b01101011000100110010: color_data = 12'b111101110000;
20'b01101011000100110011: color_data = 12'b111101110000;
20'b01101011000100110100: color_data = 12'b111101110000;
20'b01101011000100110101: color_data = 12'b111101110000;
20'b01101011000100111001: color_data = 12'b111101110000;
20'b01101011000100111010: color_data = 12'b111101110000;
20'b01101011000100111011: color_data = 12'b111101110000;
20'b01101011000100111100: color_data = 12'b111101110000;
20'b01101011000100111101: color_data = 12'b111101110000;
20'b01101011000100111110: color_data = 12'b111101110000;
20'b01101011000100111111: color_data = 12'b111101110000;
20'b01101011000101000000: color_data = 12'b111101110000;
20'b01101011000101000001: color_data = 12'b111101110000;
20'b01101011000101000010: color_data = 12'b111101110000;
20'b01101011000101000011: color_data = 12'b111101110000;
20'b01101011000101000100: color_data = 12'b111101110000;
20'b01101011000101000101: color_data = 12'b111101110000;
20'b01101011000101000110: color_data = 12'b111101110000;
20'b01101011000101000111: color_data = 12'b111101110000;
20'b01101011000101001000: color_data = 12'b111101110000;
20'b01101011000101001001: color_data = 12'b111101110000;
20'b01101011000101001010: color_data = 12'b111101110000;
20'b01101011000101001110: color_data = 12'b000011110000;
20'b01101011000101001111: color_data = 12'b000011110000;
20'b01101011000101010000: color_data = 12'b000011110000;
20'b01101011000101010001: color_data = 12'b000011110000;
20'b01101011000101010010: color_data = 12'b000011110000;
20'b01101011000101010011: color_data = 12'b000011110000;
20'b01101011000101010100: color_data = 12'b000011110000;
20'b01101011000101010101: color_data = 12'b000011110000;
20'b01101011000101010110: color_data = 12'b000011110000;
20'b01101011000101010111: color_data = 12'b000011110000;
20'b01101011000101011000: color_data = 12'b000011110000;
20'b01101011000101011001: color_data = 12'b000011110000;
20'b01101011000101011010: color_data = 12'b000011110000;
20'b01101011000101011011: color_data = 12'b000011110000;
20'b01101011000101011100: color_data = 12'b000011110000;
20'b01101011000101011101: color_data = 12'b000011110000;
20'b01101011000101011110: color_data = 12'b000011110000;
20'b01101011000101011111: color_data = 12'b000011110000;
20'b01101011000101100011: color_data = 12'b111100001111;
20'b01101011000101100100: color_data = 12'b111100001111;
20'b01101011000101100101: color_data = 12'b111100001111;
20'b01101011000101100110: color_data = 12'b111100001111;
20'b01101011000101100111: color_data = 12'b111100001111;
20'b01101011000101101000: color_data = 12'b111100001111;
20'b01101011000101101001: color_data = 12'b111100001111;
20'b01101011000101101010: color_data = 12'b111100001111;
20'b01101011000101101011: color_data = 12'b111100001111;
20'b01101011000101101100: color_data = 12'b111100001111;
20'b01101011000101101101: color_data = 12'b111100001111;
20'b01101011000101101110: color_data = 12'b111100001111;
20'b01101011000101101111: color_data = 12'b111100001111;
20'b01101011000101110000: color_data = 12'b111100001111;
20'b01101011000101110001: color_data = 12'b111100001111;
20'b01101011000101110010: color_data = 12'b111100001111;
20'b01101011000101110011: color_data = 12'b111100001111;
20'b01101011000101110100: color_data = 12'b111100001111;
20'b01101011000101111000: color_data = 12'b111100000000;
20'b01101011000101111001: color_data = 12'b111100000000;
20'b01101011000101111010: color_data = 12'b111100000000;
20'b01101011000101111011: color_data = 12'b111100000000;
20'b01101011000101111100: color_data = 12'b111100000000;
20'b01101011000101111101: color_data = 12'b111100000000;
20'b01101011000101111110: color_data = 12'b111100000000;
20'b01101011000101111111: color_data = 12'b111100000000;
20'b01101011000110000000: color_data = 12'b111100000000;
20'b01101011000110000001: color_data = 12'b111100000000;
20'b01101011000110000010: color_data = 12'b111100000000;
20'b01101011000110000011: color_data = 12'b111100000000;
20'b01101011000110000100: color_data = 12'b111100000000;
20'b01101011000110000101: color_data = 12'b111100000000;
20'b01101011000110000110: color_data = 12'b111100000000;
20'b01101011000110000111: color_data = 12'b111100000000;
20'b01101011000110001000: color_data = 12'b111100000000;
20'b01101011000110001001: color_data = 12'b111100000000;
20'b01101011000110001101: color_data = 12'b111100000000;
20'b01101011000110001110: color_data = 12'b111100000000;
20'b01101011000110001111: color_data = 12'b111100000000;
20'b01101011000110010000: color_data = 12'b111100000000;
20'b01101011000110010001: color_data = 12'b111100000000;
20'b01101011000110010010: color_data = 12'b111100000000;
20'b01101011000110010011: color_data = 12'b111100000000;
20'b01101011000110010100: color_data = 12'b111100000000;
20'b01101011000110010101: color_data = 12'b111100000000;
20'b01101011000110010110: color_data = 12'b111100000000;
20'b01101011000110010111: color_data = 12'b111100000000;
20'b01101011000110011000: color_data = 12'b111100000000;
20'b01101011000110011001: color_data = 12'b111100000000;
20'b01101011000110011010: color_data = 12'b111100000000;
20'b01101011000110011011: color_data = 12'b111100000000;
20'b01101011000110011100: color_data = 12'b111100000000;
20'b01101011000110011101: color_data = 12'b111100000000;
20'b01101011000110011110: color_data = 12'b111100000000;
20'b01101011010011111010: color_data = 12'b111101110000;
20'b01101011010011111011: color_data = 12'b111101110000;
20'b01101011010011111100: color_data = 12'b111101110000;
20'b01101011010011111101: color_data = 12'b111101110000;
20'b01101011010011111110: color_data = 12'b111101110000;
20'b01101011010011111111: color_data = 12'b111101110000;
20'b01101011010100000000: color_data = 12'b111101110000;
20'b01101011010100000001: color_data = 12'b111101110000;
20'b01101011010100000010: color_data = 12'b111101110000;
20'b01101011010100000011: color_data = 12'b111101110000;
20'b01101011010100000100: color_data = 12'b111101110000;
20'b01101011010100000101: color_data = 12'b111101110000;
20'b01101011010100000110: color_data = 12'b111101110000;
20'b01101011010100000111: color_data = 12'b111101110000;
20'b01101011010100001000: color_data = 12'b111101110000;
20'b01101011010100001001: color_data = 12'b111101110000;
20'b01101011010100001010: color_data = 12'b111101110000;
20'b01101011010100001011: color_data = 12'b111101110000;
20'b01101011010100001111: color_data = 12'b111101110000;
20'b01101011010100010000: color_data = 12'b111101110000;
20'b01101011010100010001: color_data = 12'b111101110000;
20'b01101011010100010010: color_data = 12'b111101110000;
20'b01101011010100010011: color_data = 12'b111101110000;
20'b01101011010100010100: color_data = 12'b111101110000;
20'b01101011010100010101: color_data = 12'b111101110000;
20'b01101011010100010110: color_data = 12'b111101110000;
20'b01101011010100010111: color_data = 12'b111101110000;
20'b01101011010100011000: color_data = 12'b111101110000;
20'b01101011010100011001: color_data = 12'b111101110000;
20'b01101011010100011010: color_data = 12'b111101110000;
20'b01101011010100011011: color_data = 12'b111101110000;
20'b01101011010100011100: color_data = 12'b111101110000;
20'b01101011010100011101: color_data = 12'b111101110000;
20'b01101011010100011110: color_data = 12'b111101110000;
20'b01101011010100011111: color_data = 12'b111101110000;
20'b01101011010100100000: color_data = 12'b111101110000;
20'b01101011010100100100: color_data = 12'b111101110000;
20'b01101011010100100101: color_data = 12'b111101110000;
20'b01101011010100100110: color_data = 12'b111101110000;
20'b01101011010100100111: color_data = 12'b111101110000;
20'b01101011010100101000: color_data = 12'b111101110000;
20'b01101011010100101001: color_data = 12'b111101110000;
20'b01101011010100101010: color_data = 12'b111101110000;
20'b01101011010100101011: color_data = 12'b111101110000;
20'b01101011010100101100: color_data = 12'b111101110000;
20'b01101011010100101101: color_data = 12'b111101110000;
20'b01101011010100101110: color_data = 12'b111101110000;
20'b01101011010100101111: color_data = 12'b111101110000;
20'b01101011010100110000: color_data = 12'b111101110000;
20'b01101011010100110001: color_data = 12'b111101110000;
20'b01101011010100110010: color_data = 12'b111101110000;
20'b01101011010100110011: color_data = 12'b111101110000;
20'b01101011010100110100: color_data = 12'b111101110000;
20'b01101011010100110101: color_data = 12'b111101110000;
20'b01101011010100111001: color_data = 12'b111101110000;
20'b01101011010100111010: color_data = 12'b111101110000;
20'b01101011010100111011: color_data = 12'b111101110000;
20'b01101011010100111100: color_data = 12'b111101110000;
20'b01101011010100111101: color_data = 12'b111101110000;
20'b01101011010100111110: color_data = 12'b111101110000;
20'b01101011010100111111: color_data = 12'b111101110000;
20'b01101011010101000000: color_data = 12'b111101110000;
20'b01101011010101000001: color_data = 12'b111101110000;
20'b01101011010101000010: color_data = 12'b111101110000;
20'b01101011010101000011: color_data = 12'b111101110000;
20'b01101011010101000100: color_data = 12'b111101110000;
20'b01101011010101000101: color_data = 12'b111101110000;
20'b01101011010101000110: color_data = 12'b111101110000;
20'b01101011010101000111: color_data = 12'b111101110000;
20'b01101011010101001000: color_data = 12'b111101110000;
20'b01101011010101001001: color_data = 12'b111101110000;
20'b01101011010101001010: color_data = 12'b111101110000;
20'b01101011010101001110: color_data = 12'b000011110000;
20'b01101011010101001111: color_data = 12'b000011110000;
20'b01101011010101010000: color_data = 12'b000011110000;
20'b01101011010101010001: color_data = 12'b000011110000;
20'b01101011010101010010: color_data = 12'b000011110000;
20'b01101011010101010011: color_data = 12'b000011110000;
20'b01101011010101010100: color_data = 12'b000011110000;
20'b01101011010101010101: color_data = 12'b000011110000;
20'b01101011010101010110: color_data = 12'b000011110000;
20'b01101011010101010111: color_data = 12'b000011110000;
20'b01101011010101011000: color_data = 12'b000011110000;
20'b01101011010101011001: color_data = 12'b000011110000;
20'b01101011010101011010: color_data = 12'b000011110000;
20'b01101011010101011011: color_data = 12'b000011110000;
20'b01101011010101011100: color_data = 12'b000011110000;
20'b01101011010101011101: color_data = 12'b000011110000;
20'b01101011010101011110: color_data = 12'b000011110000;
20'b01101011010101011111: color_data = 12'b000011110000;
20'b01101011010101100011: color_data = 12'b111100001111;
20'b01101011010101100100: color_data = 12'b111100001111;
20'b01101011010101100101: color_data = 12'b111100001111;
20'b01101011010101100110: color_data = 12'b111100001111;
20'b01101011010101100111: color_data = 12'b111100001111;
20'b01101011010101101000: color_data = 12'b111100001111;
20'b01101011010101101001: color_data = 12'b111100001111;
20'b01101011010101101010: color_data = 12'b111100001111;
20'b01101011010101101011: color_data = 12'b111100001111;
20'b01101011010101101100: color_data = 12'b111100001111;
20'b01101011010101101101: color_data = 12'b111100001111;
20'b01101011010101101110: color_data = 12'b111100001111;
20'b01101011010101101111: color_data = 12'b111100001111;
20'b01101011010101110000: color_data = 12'b111100001111;
20'b01101011010101110001: color_data = 12'b111100001111;
20'b01101011010101110010: color_data = 12'b111100001111;
20'b01101011010101110011: color_data = 12'b111100001111;
20'b01101011010101110100: color_data = 12'b111100001111;
20'b01101011010101111000: color_data = 12'b111100000000;
20'b01101011010101111001: color_data = 12'b111100000000;
20'b01101011010101111010: color_data = 12'b111100000000;
20'b01101011010101111011: color_data = 12'b111100000000;
20'b01101011010101111100: color_data = 12'b111100000000;
20'b01101011010101111101: color_data = 12'b111100000000;
20'b01101011010101111110: color_data = 12'b111100000000;
20'b01101011010101111111: color_data = 12'b111100000000;
20'b01101011010110000000: color_data = 12'b111100000000;
20'b01101011010110000001: color_data = 12'b111100000000;
20'b01101011010110000010: color_data = 12'b111100000000;
20'b01101011010110000011: color_data = 12'b111100000000;
20'b01101011010110000100: color_data = 12'b111100000000;
20'b01101011010110000101: color_data = 12'b111100000000;
20'b01101011010110000110: color_data = 12'b111100000000;
20'b01101011010110000111: color_data = 12'b111100000000;
20'b01101011010110001000: color_data = 12'b111100000000;
20'b01101011010110001001: color_data = 12'b111100000000;
20'b01101011010110001101: color_data = 12'b111100000000;
20'b01101011010110001110: color_data = 12'b111100000000;
20'b01101011010110001111: color_data = 12'b111100000000;
20'b01101011010110010000: color_data = 12'b111100000000;
20'b01101011010110010001: color_data = 12'b111100000000;
20'b01101011010110010010: color_data = 12'b111100000000;
20'b01101011010110010011: color_data = 12'b111100000000;
20'b01101011010110010100: color_data = 12'b111100000000;
20'b01101011010110010101: color_data = 12'b111100000000;
20'b01101011010110010110: color_data = 12'b111100000000;
20'b01101011010110010111: color_data = 12'b111100000000;
20'b01101011010110011000: color_data = 12'b111100000000;
20'b01101011010110011001: color_data = 12'b111100000000;
20'b01101011010110011010: color_data = 12'b111100000000;
20'b01101011010110011011: color_data = 12'b111100000000;
20'b01101011010110011100: color_data = 12'b111100000000;
20'b01101011010110011101: color_data = 12'b111100000000;
20'b01101011010110011110: color_data = 12'b111100000000;
20'b01101011100011111010: color_data = 12'b111101110000;
20'b01101011100011111011: color_data = 12'b111101110000;
20'b01101011100011111100: color_data = 12'b111101110000;
20'b01101011100011111101: color_data = 12'b111101110000;
20'b01101011100011111110: color_data = 12'b111101110000;
20'b01101011100011111111: color_data = 12'b111101110000;
20'b01101011100100000000: color_data = 12'b111101110000;
20'b01101011100100000001: color_data = 12'b111101110000;
20'b01101011100100000010: color_data = 12'b111101110000;
20'b01101011100100000011: color_data = 12'b111101110000;
20'b01101011100100000100: color_data = 12'b111101110000;
20'b01101011100100000101: color_data = 12'b111101110000;
20'b01101011100100000110: color_data = 12'b111101110000;
20'b01101011100100000111: color_data = 12'b111101110000;
20'b01101011100100001000: color_data = 12'b111101110000;
20'b01101011100100001001: color_data = 12'b111101110000;
20'b01101011100100001010: color_data = 12'b111101110000;
20'b01101011100100001011: color_data = 12'b111101110000;
20'b01101011100100001111: color_data = 12'b111101110000;
20'b01101011100100010000: color_data = 12'b111101110000;
20'b01101011100100010001: color_data = 12'b111101110000;
20'b01101011100100010010: color_data = 12'b111101110000;
20'b01101011100100010011: color_data = 12'b111101110000;
20'b01101011100100010100: color_data = 12'b111101110000;
20'b01101011100100010101: color_data = 12'b111101110000;
20'b01101011100100010110: color_data = 12'b111101110000;
20'b01101011100100010111: color_data = 12'b111101110000;
20'b01101011100100011000: color_data = 12'b111101110000;
20'b01101011100100011001: color_data = 12'b111101110000;
20'b01101011100100011010: color_data = 12'b111101110000;
20'b01101011100100011011: color_data = 12'b111101110000;
20'b01101011100100011100: color_data = 12'b111101110000;
20'b01101011100100011101: color_data = 12'b111101110000;
20'b01101011100100011110: color_data = 12'b111101110000;
20'b01101011100100011111: color_data = 12'b111101110000;
20'b01101011100100100000: color_data = 12'b111101110000;
20'b01101011100100100100: color_data = 12'b111101110000;
20'b01101011100100100101: color_data = 12'b111101110000;
20'b01101011100100100110: color_data = 12'b111101110000;
20'b01101011100100100111: color_data = 12'b111101110000;
20'b01101011100100101000: color_data = 12'b111101110000;
20'b01101011100100101001: color_data = 12'b111101110000;
20'b01101011100100101010: color_data = 12'b111101110000;
20'b01101011100100101011: color_data = 12'b111101110000;
20'b01101011100100101100: color_data = 12'b111101110000;
20'b01101011100100101101: color_data = 12'b111101110000;
20'b01101011100100101110: color_data = 12'b111101110000;
20'b01101011100100101111: color_data = 12'b111101110000;
20'b01101011100100110000: color_data = 12'b111101110000;
20'b01101011100100110001: color_data = 12'b111101110000;
20'b01101011100100110010: color_data = 12'b111101110000;
20'b01101011100100110011: color_data = 12'b111101110000;
20'b01101011100100110100: color_data = 12'b111101110000;
20'b01101011100100110101: color_data = 12'b111101110000;
20'b01101011100100111001: color_data = 12'b111101110000;
20'b01101011100100111010: color_data = 12'b111101110000;
20'b01101011100100111011: color_data = 12'b111101110000;
20'b01101011100100111100: color_data = 12'b111101110000;
20'b01101011100100111101: color_data = 12'b111101110000;
20'b01101011100100111110: color_data = 12'b111101110000;
20'b01101011100100111111: color_data = 12'b111101110000;
20'b01101011100101000000: color_data = 12'b111101110000;
20'b01101011100101000001: color_data = 12'b111101110000;
20'b01101011100101000010: color_data = 12'b111101110000;
20'b01101011100101000011: color_data = 12'b111101110000;
20'b01101011100101000100: color_data = 12'b111101110000;
20'b01101011100101000101: color_data = 12'b111101110000;
20'b01101011100101000110: color_data = 12'b111101110000;
20'b01101011100101000111: color_data = 12'b111101110000;
20'b01101011100101001000: color_data = 12'b111101110000;
20'b01101011100101001001: color_data = 12'b111101110000;
20'b01101011100101001010: color_data = 12'b111101110000;
20'b01101011100101001110: color_data = 12'b000011110000;
20'b01101011100101001111: color_data = 12'b000011110000;
20'b01101011100101010000: color_data = 12'b000011110000;
20'b01101011100101010001: color_data = 12'b000011110000;
20'b01101011100101010010: color_data = 12'b000011110000;
20'b01101011100101010011: color_data = 12'b000011110000;
20'b01101011100101010100: color_data = 12'b000011110000;
20'b01101011100101010101: color_data = 12'b000011110000;
20'b01101011100101010110: color_data = 12'b000011110000;
20'b01101011100101010111: color_data = 12'b000011110000;
20'b01101011100101011000: color_data = 12'b000011110000;
20'b01101011100101011001: color_data = 12'b000011110000;
20'b01101011100101011010: color_data = 12'b000011110000;
20'b01101011100101011011: color_data = 12'b000011110000;
20'b01101011100101011100: color_data = 12'b000011110000;
20'b01101011100101011101: color_data = 12'b000011110000;
20'b01101011100101011110: color_data = 12'b000011110000;
20'b01101011100101011111: color_data = 12'b000011110000;
20'b01101011100101100011: color_data = 12'b111100001111;
20'b01101011100101100100: color_data = 12'b111100001111;
20'b01101011100101100101: color_data = 12'b111100001111;
20'b01101011100101100110: color_data = 12'b111100001111;
20'b01101011100101100111: color_data = 12'b111100001111;
20'b01101011100101101000: color_data = 12'b111100001111;
20'b01101011100101101001: color_data = 12'b111100001111;
20'b01101011100101101010: color_data = 12'b111100001111;
20'b01101011100101101011: color_data = 12'b111100001111;
20'b01101011100101101100: color_data = 12'b111100001111;
20'b01101011100101101101: color_data = 12'b111100001111;
20'b01101011100101101110: color_data = 12'b111100001111;
20'b01101011100101101111: color_data = 12'b111100001111;
20'b01101011100101110000: color_data = 12'b111100001111;
20'b01101011100101110001: color_data = 12'b111100001111;
20'b01101011100101110010: color_data = 12'b111100001111;
20'b01101011100101110011: color_data = 12'b111100001111;
20'b01101011100101110100: color_data = 12'b111100001111;
20'b01101011100101111000: color_data = 12'b111100000000;
20'b01101011100101111001: color_data = 12'b111100000000;
20'b01101011100101111010: color_data = 12'b111100000000;
20'b01101011100101111011: color_data = 12'b111100000000;
20'b01101011100101111100: color_data = 12'b111100000000;
20'b01101011100101111101: color_data = 12'b111100000000;
20'b01101011100101111110: color_data = 12'b111100000000;
20'b01101011100101111111: color_data = 12'b111100000000;
20'b01101011100110000000: color_data = 12'b111100000000;
20'b01101011100110000001: color_data = 12'b111100000000;
20'b01101011100110000010: color_data = 12'b111100000000;
20'b01101011100110000011: color_data = 12'b111100000000;
20'b01101011100110000100: color_data = 12'b111100000000;
20'b01101011100110000101: color_data = 12'b111100000000;
20'b01101011100110000110: color_data = 12'b111100000000;
20'b01101011100110000111: color_data = 12'b111100000000;
20'b01101011100110001000: color_data = 12'b111100000000;
20'b01101011100110001001: color_data = 12'b111100000000;
20'b01101011100110001101: color_data = 12'b111100000000;
20'b01101011100110001110: color_data = 12'b111100000000;
20'b01101011100110001111: color_data = 12'b111100000000;
20'b01101011100110010000: color_data = 12'b111100000000;
20'b01101011100110010001: color_data = 12'b111100000000;
20'b01101011100110010010: color_data = 12'b111100000000;
20'b01101011100110010011: color_data = 12'b111100000000;
20'b01101011100110010100: color_data = 12'b111100000000;
20'b01101011100110010101: color_data = 12'b111100000000;
20'b01101011100110010110: color_data = 12'b111100000000;
20'b01101011100110010111: color_data = 12'b111100000000;
20'b01101011100110011000: color_data = 12'b111100000000;
20'b01101011100110011001: color_data = 12'b111100000000;
20'b01101011100110011010: color_data = 12'b111100000000;
20'b01101011100110011011: color_data = 12'b111100000000;
20'b01101011100110011100: color_data = 12'b111100000000;
20'b01101011100110011101: color_data = 12'b111100000000;
20'b01101011100110011110: color_data = 12'b111100000000;
20'b01101011110011111010: color_data = 12'b111101110000;
20'b01101011110011111011: color_data = 12'b111101110000;
20'b01101011110011111100: color_data = 12'b111101110000;
20'b01101011110011111101: color_data = 12'b111101110000;
20'b01101011110011111110: color_data = 12'b111101110000;
20'b01101011110011111111: color_data = 12'b111101110000;
20'b01101011110100000000: color_data = 12'b111101110000;
20'b01101011110100000001: color_data = 12'b111101110000;
20'b01101011110100000010: color_data = 12'b111101110000;
20'b01101011110100000011: color_data = 12'b111101110000;
20'b01101011110100000100: color_data = 12'b111101110000;
20'b01101011110100000101: color_data = 12'b111101110000;
20'b01101011110100000110: color_data = 12'b111101110000;
20'b01101011110100000111: color_data = 12'b111101110000;
20'b01101011110100001000: color_data = 12'b111101110000;
20'b01101011110100001001: color_data = 12'b111101110000;
20'b01101011110100001010: color_data = 12'b111101110000;
20'b01101011110100001011: color_data = 12'b111101110000;
20'b01101011110100001111: color_data = 12'b111101110000;
20'b01101011110100010000: color_data = 12'b111101110000;
20'b01101011110100010001: color_data = 12'b111101110000;
20'b01101011110100010010: color_data = 12'b111101110000;
20'b01101011110100010011: color_data = 12'b111101110000;
20'b01101011110100010100: color_data = 12'b111101110000;
20'b01101011110100010101: color_data = 12'b111101110000;
20'b01101011110100010110: color_data = 12'b111101110000;
20'b01101011110100010111: color_data = 12'b111101110000;
20'b01101011110100011000: color_data = 12'b111101110000;
20'b01101011110100011001: color_data = 12'b111101110000;
20'b01101011110100011010: color_data = 12'b111101110000;
20'b01101011110100011011: color_data = 12'b111101110000;
20'b01101011110100011100: color_data = 12'b111101110000;
20'b01101011110100011101: color_data = 12'b111101110000;
20'b01101011110100011110: color_data = 12'b111101110000;
20'b01101011110100011111: color_data = 12'b111101110000;
20'b01101011110100100000: color_data = 12'b111101110000;
20'b01101011110100100100: color_data = 12'b111101110000;
20'b01101011110100100101: color_data = 12'b111101110000;
20'b01101011110100100110: color_data = 12'b111101110000;
20'b01101011110100100111: color_data = 12'b111101110000;
20'b01101011110100101000: color_data = 12'b111101110000;
20'b01101011110100101001: color_data = 12'b111101110000;
20'b01101011110100101010: color_data = 12'b111101110000;
20'b01101011110100101011: color_data = 12'b111101110000;
20'b01101011110100101100: color_data = 12'b111101110000;
20'b01101011110100101101: color_data = 12'b111101110000;
20'b01101011110100101110: color_data = 12'b111101110000;
20'b01101011110100101111: color_data = 12'b111101110000;
20'b01101011110100110000: color_data = 12'b111101110000;
20'b01101011110100110001: color_data = 12'b111101110000;
20'b01101011110100110010: color_data = 12'b111101110000;
20'b01101011110100110011: color_data = 12'b111101110000;
20'b01101011110100110100: color_data = 12'b111101110000;
20'b01101011110100110101: color_data = 12'b111101110000;
20'b01101011110100111001: color_data = 12'b111101110000;
20'b01101011110100111010: color_data = 12'b111101110000;
20'b01101011110100111011: color_data = 12'b111101110000;
20'b01101011110100111100: color_data = 12'b111101110000;
20'b01101011110100111101: color_data = 12'b111101110000;
20'b01101011110100111110: color_data = 12'b111101110000;
20'b01101011110100111111: color_data = 12'b111101110000;
20'b01101011110101000000: color_data = 12'b111101110000;
20'b01101011110101000001: color_data = 12'b111101110000;
20'b01101011110101000010: color_data = 12'b111101110000;
20'b01101011110101000011: color_data = 12'b111101110000;
20'b01101011110101000100: color_data = 12'b111101110000;
20'b01101011110101000101: color_data = 12'b111101110000;
20'b01101011110101000110: color_data = 12'b111101110000;
20'b01101011110101000111: color_data = 12'b111101110000;
20'b01101011110101001000: color_data = 12'b111101110000;
20'b01101011110101001001: color_data = 12'b111101110000;
20'b01101011110101001010: color_data = 12'b111101110000;
20'b01101011110101001110: color_data = 12'b000011110000;
20'b01101011110101001111: color_data = 12'b000011110000;
20'b01101011110101010000: color_data = 12'b000011110000;
20'b01101011110101010001: color_data = 12'b000011110000;
20'b01101011110101010010: color_data = 12'b000011110000;
20'b01101011110101010011: color_data = 12'b000011110000;
20'b01101011110101010100: color_data = 12'b000011110000;
20'b01101011110101010101: color_data = 12'b000011110000;
20'b01101011110101010110: color_data = 12'b000011110000;
20'b01101011110101010111: color_data = 12'b000011110000;
20'b01101011110101011000: color_data = 12'b000011110000;
20'b01101011110101011001: color_data = 12'b000011110000;
20'b01101011110101011010: color_data = 12'b000011110000;
20'b01101011110101011011: color_data = 12'b000011110000;
20'b01101011110101011100: color_data = 12'b000011110000;
20'b01101011110101011101: color_data = 12'b000011110000;
20'b01101011110101011110: color_data = 12'b000011110000;
20'b01101011110101011111: color_data = 12'b000011110000;
20'b01101011110101100011: color_data = 12'b111100001111;
20'b01101011110101100100: color_data = 12'b111100001111;
20'b01101011110101100101: color_data = 12'b111100001111;
20'b01101011110101100110: color_data = 12'b111100001111;
20'b01101011110101100111: color_data = 12'b111100001111;
20'b01101011110101101000: color_data = 12'b111100001111;
20'b01101011110101101001: color_data = 12'b111100001111;
20'b01101011110101101010: color_data = 12'b111100001111;
20'b01101011110101101011: color_data = 12'b111100001111;
20'b01101011110101101100: color_data = 12'b111100001111;
20'b01101011110101101101: color_data = 12'b111100001111;
20'b01101011110101101110: color_data = 12'b111100001111;
20'b01101011110101101111: color_data = 12'b111100001111;
20'b01101011110101110000: color_data = 12'b111100001111;
20'b01101011110101110001: color_data = 12'b111100001111;
20'b01101011110101110010: color_data = 12'b111100001111;
20'b01101011110101110011: color_data = 12'b111100001111;
20'b01101011110101110100: color_data = 12'b111100001111;
20'b01101011110101111000: color_data = 12'b111100000000;
20'b01101011110101111001: color_data = 12'b111100000000;
20'b01101011110101111010: color_data = 12'b111100000000;
20'b01101011110101111011: color_data = 12'b111100000000;
20'b01101011110101111100: color_data = 12'b111100000000;
20'b01101011110101111101: color_data = 12'b111100000000;
20'b01101011110101111110: color_data = 12'b111100000000;
20'b01101011110101111111: color_data = 12'b111100000000;
20'b01101011110110000000: color_data = 12'b111100000000;
20'b01101011110110000001: color_data = 12'b111100000000;
20'b01101011110110000010: color_data = 12'b111100000000;
20'b01101011110110000011: color_data = 12'b111100000000;
20'b01101011110110000100: color_data = 12'b111100000000;
20'b01101011110110000101: color_data = 12'b111100000000;
20'b01101011110110000110: color_data = 12'b111100000000;
20'b01101011110110000111: color_data = 12'b111100000000;
20'b01101011110110001000: color_data = 12'b111100000000;
20'b01101011110110001001: color_data = 12'b111100000000;
20'b01101011110110001101: color_data = 12'b111100000000;
20'b01101011110110001110: color_data = 12'b111100000000;
20'b01101011110110001111: color_data = 12'b111100000000;
20'b01101011110110010000: color_data = 12'b111100000000;
20'b01101011110110010001: color_data = 12'b111100000000;
20'b01101011110110010010: color_data = 12'b111100000000;
20'b01101011110110010011: color_data = 12'b111100000000;
20'b01101011110110010100: color_data = 12'b111100000000;
20'b01101011110110010101: color_data = 12'b111100000000;
20'b01101011110110010110: color_data = 12'b111100000000;
20'b01101011110110010111: color_data = 12'b111100000000;
20'b01101011110110011000: color_data = 12'b111100000000;
20'b01101011110110011001: color_data = 12'b111100000000;
20'b01101011110110011010: color_data = 12'b111100000000;
20'b01101011110110011011: color_data = 12'b111100000000;
20'b01101011110110011100: color_data = 12'b111100000000;
20'b01101011110110011101: color_data = 12'b111100000000;
20'b01101011110110011110: color_data = 12'b111100000000;
20'b01101100000011111010: color_data = 12'b111101110000;
20'b01101100000011111011: color_data = 12'b111101110000;
20'b01101100000011111100: color_data = 12'b111101110000;
20'b01101100000011111101: color_data = 12'b111101110000;
20'b01101100000011111110: color_data = 12'b111101110000;
20'b01101100000011111111: color_data = 12'b111101110000;
20'b01101100000100000000: color_data = 12'b111101110000;
20'b01101100000100000001: color_data = 12'b111101110000;
20'b01101100000100000010: color_data = 12'b111101110000;
20'b01101100000100000011: color_data = 12'b111101110000;
20'b01101100000100000100: color_data = 12'b111101110000;
20'b01101100000100000101: color_data = 12'b111101110000;
20'b01101100000100000110: color_data = 12'b111101110000;
20'b01101100000100000111: color_data = 12'b111101110000;
20'b01101100000100001000: color_data = 12'b111101110000;
20'b01101100000100001001: color_data = 12'b111101110000;
20'b01101100000100001010: color_data = 12'b111101110000;
20'b01101100000100001011: color_data = 12'b111101110000;
20'b01101100000100001111: color_data = 12'b111101110000;
20'b01101100000100010000: color_data = 12'b111101110000;
20'b01101100000100010001: color_data = 12'b111101110000;
20'b01101100000100010010: color_data = 12'b111101110000;
20'b01101100000100010011: color_data = 12'b111101110000;
20'b01101100000100010100: color_data = 12'b111101110000;
20'b01101100000100010101: color_data = 12'b111101110000;
20'b01101100000100010110: color_data = 12'b111101110000;
20'b01101100000100010111: color_data = 12'b111101110000;
20'b01101100000100011000: color_data = 12'b111101110000;
20'b01101100000100011001: color_data = 12'b111101110000;
20'b01101100000100011010: color_data = 12'b111101110000;
20'b01101100000100011011: color_data = 12'b111101110000;
20'b01101100000100011100: color_data = 12'b111101110000;
20'b01101100000100011101: color_data = 12'b111101110000;
20'b01101100000100011110: color_data = 12'b111101110000;
20'b01101100000100011111: color_data = 12'b111101110000;
20'b01101100000100100000: color_data = 12'b111101110000;
20'b01101100000100100100: color_data = 12'b111101110000;
20'b01101100000100100101: color_data = 12'b111101110000;
20'b01101100000100100110: color_data = 12'b111101110000;
20'b01101100000100100111: color_data = 12'b111101110000;
20'b01101100000100101000: color_data = 12'b111101110000;
20'b01101100000100101001: color_data = 12'b111101110000;
20'b01101100000100101010: color_data = 12'b111101110000;
20'b01101100000100101011: color_data = 12'b111101110000;
20'b01101100000100101100: color_data = 12'b111101110000;
20'b01101100000100101101: color_data = 12'b111101110000;
20'b01101100000100101110: color_data = 12'b111101110000;
20'b01101100000100101111: color_data = 12'b111101110000;
20'b01101100000100110000: color_data = 12'b111101110000;
20'b01101100000100110001: color_data = 12'b111101110000;
20'b01101100000100110010: color_data = 12'b111101110000;
20'b01101100000100110011: color_data = 12'b111101110000;
20'b01101100000100110100: color_data = 12'b111101110000;
20'b01101100000100110101: color_data = 12'b111101110000;
20'b01101100000100111001: color_data = 12'b111101110000;
20'b01101100000100111010: color_data = 12'b111101110000;
20'b01101100000100111011: color_data = 12'b111101110000;
20'b01101100000100111100: color_data = 12'b111101110000;
20'b01101100000100111101: color_data = 12'b111101110000;
20'b01101100000100111110: color_data = 12'b111101110000;
20'b01101100000100111111: color_data = 12'b111101110000;
20'b01101100000101000000: color_data = 12'b111101110000;
20'b01101100000101000001: color_data = 12'b111101110000;
20'b01101100000101000010: color_data = 12'b111101110000;
20'b01101100000101000011: color_data = 12'b111101110000;
20'b01101100000101000100: color_data = 12'b111101110000;
20'b01101100000101000101: color_data = 12'b111101110000;
20'b01101100000101000110: color_data = 12'b111101110000;
20'b01101100000101000111: color_data = 12'b111101110000;
20'b01101100000101001000: color_data = 12'b111101110000;
20'b01101100000101001001: color_data = 12'b111101110000;
20'b01101100000101001010: color_data = 12'b111101110000;
20'b01101100000101001110: color_data = 12'b000011110000;
20'b01101100000101001111: color_data = 12'b000011110000;
20'b01101100000101010000: color_data = 12'b000011110000;
20'b01101100000101010001: color_data = 12'b000011110000;
20'b01101100000101010010: color_data = 12'b000011110000;
20'b01101100000101010011: color_data = 12'b000011110000;
20'b01101100000101010100: color_data = 12'b000011110000;
20'b01101100000101010101: color_data = 12'b000011110000;
20'b01101100000101010110: color_data = 12'b000011110000;
20'b01101100000101010111: color_data = 12'b000011110000;
20'b01101100000101011000: color_data = 12'b000011110000;
20'b01101100000101011001: color_data = 12'b000011110000;
20'b01101100000101011010: color_data = 12'b000011110000;
20'b01101100000101011011: color_data = 12'b000011110000;
20'b01101100000101011100: color_data = 12'b000011110000;
20'b01101100000101011101: color_data = 12'b000011110000;
20'b01101100000101011110: color_data = 12'b000011110000;
20'b01101100000101011111: color_data = 12'b000011110000;
20'b01101100000101100011: color_data = 12'b111100001111;
20'b01101100000101100100: color_data = 12'b111100001111;
20'b01101100000101100101: color_data = 12'b111100001111;
20'b01101100000101100110: color_data = 12'b111100001111;
20'b01101100000101100111: color_data = 12'b111100001111;
20'b01101100000101101000: color_data = 12'b111100001111;
20'b01101100000101101001: color_data = 12'b111100001111;
20'b01101100000101101010: color_data = 12'b111100001111;
20'b01101100000101101011: color_data = 12'b111100001111;
20'b01101100000101101100: color_data = 12'b111100001111;
20'b01101100000101101101: color_data = 12'b111100001111;
20'b01101100000101101110: color_data = 12'b111100001111;
20'b01101100000101101111: color_data = 12'b111100001111;
20'b01101100000101110000: color_data = 12'b111100001111;
20'b01101100000101110001: color_data = 12'b111100001111;
20'b01101100000101110010: color_data = 12'b111100001111;
20'b01101100000101110011: color_data = 12'b111100001111;
20'b01101100000101110100: color_data = 12'b111100001111;
20'b01101100000101111000: color_data = 12'b111100000000;
20'b01101100000101111001: color_data = 12'b111100000000;
20'b01101100000101111010: color_data = 12'b111100000000;
20'b01101100000101111011: color_data = 12'b111100000000;
20'b01101100000101111100: color_data = 12'b111100000000;
20'b01101100000101111101: color_data = 12'b111100000000;
20'b01101100000101111110: color_data = 12'b111100000000;
20'b01101100000101111111: color_data = 12'b111100000000;
20'b01101100000110000000: color_data = 12'b111100000000;
20'b01101100000110000001: color_data = 12'b111100000000;
20'b01101100000110000010: color_data = 12'b111100000000;
20'b01101100000110000011: color_data = 12'b111100000000;
20'b01101100000110000100: color_data = 12'b111100000000;
20'b01101100000110000101: color_data = 12'b111100000000;
20'b01101100000110000110: color_data = 12'b111100000000;
20'b01101100000110000111: color_data = 12'b111100000000;
20'b01101100000110001000: color_data = 12'b111100000000;
20'b01101100000110001001: color_data = 12'b111100000000;
20'b01101100000110001101: color_data = 12'b111100000000;
20'b01101100000110001110: color_data = 12'b111100000000;
20'b01101100000110001111: color_data = 12'b111100000000;
20'b01101100000110010000: color_data = 12'b111100000000;
20'b01101100000110010001: color_data = 12'b111100000000;
20'b01101100000110010010: color_data = 12'b111100000000;
20'b01101100000110010011: color_data = 12'b111100000000;
20'b01101100000110010100: color_data = 12'b111100000000;
20'b01101100000110010101: color_data = 12'b111100000000;
20'b01101100000110010110: color_data = 12'b111100000000;
20'b01101100000110010111: color_data = 12'b111100000000;
20'b01101100000110011000: color_data = 12'b111100000000;
20'b01101100000110011001: color_data = 12'b111100000000;
20'b01101100000110011010: color_data = 12'b111100000000;
20'b01101100000110011011: color_data = 12'b111100000000;
20'b01101100000110011100: color_data = 12'b111100000000;
20'b01101100000110011101: color_data = 12'b111100000000;
20'b01101100000110011110: color_data = 12'b111100000000;
20'b01101100010011111010: color_data = 12'b111101110000;
20'b01101100010011111011: color_data = 12'b111101110000;
20'b01101100010011111100: color_data = 12'b111101110000;
20'b01101100010011111101: color_data = 12'b111101110000;
20'b01101100010011111110: color_data = 12'b111101110000;
20'b01101100010011111111: color_data = 12'b111101110000;
20'b01101100010100000000: color_data = 12'b111101110000;
20'b01101100010100000001: color_data = 12'b111101110000;
20'b01101100010100000010: color_data = 12'b111101110000;
20'b01101100010100000011: color_data = 12'b111101110000;
20'b01101100010100000100: color_data = 12'b111101110000;
20'b01101100010100000101: color_data = 12'b111101110000;
20'b01101100010100000110: color_data = 12'b111101110000;
20'b01101100010100000111: color_data = 12'b111101110000;
20'b01101100010100001000: color_data = 12'b111101110000;
20'b01101100010100001001: color_data = 12'b111101110000;
20'b01101100010100001010: color_data = 12'b111101110000;
20'b01101100010100001011: color_data = 12'b111101110000;
20'b01101100010100001111: color_data = 12'b111101110000;
20'b01101100010100010000: color_data = 12'b111101110000;
20'b01101100010100010001: color_data = 12'b111101110000;
20'b01101100010100010010: color_data = 12'b111101110000;
20'b01101100010100010011: color_data = 12'b111101110000;
20'b01101100010100010100: color_data = 12'b111101110000;
20'b01101100010100010101: color_data = 12'b111101110000;
20'b01101100010100010110: color_data = 12'b111101110000;
20'b01101100010100010111: color_data = 12'b111101110000;
20'b01101100010100011000: color_data = 12'b111101110000;
20'b01101100010100011001: color_data = 12'b111101110000;
20'b01101100010100011010: color_data = 12'b111101110000;
20'b01101100010100011011: color_data = 12'b111101110000;
20'b01101100010100011100: color_data = 12'b111101110000;
20'b01101100010100011101: color_data = 12'b111101110000;
20'b01101100010100011110: color_data = 12'b111101110000;
20'b01101100010100011111: color_data = 12'b111101110000;
20'b01101100010100100000: color_data = 12'b111101110000;
20'b01101100010100100100: color_data = 12'b111101110000;
20'b01101100010100100101: color_data = 12'b111101110000;
20'b01101100010100100110: color_data = 12'b111101110000;
20'b01101100010100100111: color_data = 12'b111101110000;
20'b01101100010100101000: color_data = 12'b111101110000;
20'b01101100010100101001: color_data = 12'b111101110000;
20'b01101100010100101010: color_data = 12'b111101110000;
20'b01101100010100101011: color_data = 12'b111101110000;
20'b01101100010100101100: color_data = 12'b111101110000;
20'b01101100010100101101: color_data = 12'b111101110000;
20'b01101100010100101110: color_data = 12'b111101110000;
20'b01101100010100101111: color_data = 12'b111101110000;
20'b01101100010100110000: color_data = 12'b111101110000;
20'b01101100010100110001: color_data = 12'b111101110000;
20'b01101100010100110010: color_data = 12'b111101110000;
20'b01101100010100110011: color_data = 12'b111101110000;
20'b01101100010100110100: color_data = 12'b111101110000;
20'b01101100010100110101: color_data = 12'b111101110000;
20'b01101100010100111001: color_data = 12'b111101110000;
20'b01101100010100111010: color_data = 12'b111101110000;
20'b01101100010100111011: color_data = 12'b111101110000;
20'b01101100010100111100: color_data = 12'b111101110000;
20'b01101100010100111101: color_data = 12'b111101110000;
20'b01101100010100111110: color_data = 12'b111101110000;
20'b01101100010100111111: color_data = 12'b111101110000;
20'b01101100010101000000: color_data = 12'b111101110000;
20'b01101100010101000001: color_data = 12'b111101110000;
20'b01101100010101000010: color_data = 12'b111101110000;
20'b01101100010101000011: color_data = 12'b111101110000;
20'b01101100010101000100: color_data = 12'b111101110000;
20'b01101100010101000101: color_data = 12'b111101110000;
20'b01101100010101000110: color_data = 12'b111101110000;
20'b01101100010101000111: color_data = 12'b111101110000;
20'b01101100010101001000: color_data = 12'b111101110000;
20'b01101100010101001001: color_data = 12'b111101110000;
20'b01101100010101001010: color_data = 12'b111101110000;
20'b01101100010101001110: color_data = 12'b000011110000;
20'b01101100010101001111: color_data = 12'b000011110000;
20'b01101100010101010000: color_data = 12'b000011110000;
20'b01101100010101010001: color_data = 12'b000011110000;
20'b01101100010101010010: color_data = 12'b000011110000;
20'b01101100010101010011: color_data = 12'b000011110000;
20'b01101100010101010100: color_data = 12'b000011110000;
20'b01101100010101010101: color_data = 12'b000011110000;
20'b01101100010101010110: color_data = 12'b000011110000;
20'b01101100010101010111: color_data = 12'b000011110000;
20'b01101100010101011000: color_data = 12'b000011110000;
20'b01101100010101011001: color_data = 12'b000011110000;
20'b01101100010101011010: color_data = 12'b000011110000;
20'b01101100010101011011: color_data = 12'b000011110000;
20'b01101100010101011100: color_data = 12'b000011110000;
20'b01101100010101011101: color_data = 12'b000011110000;
20'b01101100010101011110: color_data = 12'b000011110000;
20'b01101100010101011111: color_data = 12'b000011110000;
20'b01101100010101100011: color_data = 12'b111100001111;
20'b01101100010101100100: color_data = 12'b111100001111;
20'b01101100010101100101: color_data = 12'b111100001111;
20'b01101100010101100110: color_data = 12'b111100001111;
20'b01101100010101100111: color_data = 12'b111100001111;
20'b01101100010101101000: color_data = 12'b111100001111;
20'b01101100010101101001: color_data = 12'b111100001111;
20'b01101100010101101010: color_data = 12'b111100001111;
20'b01101100010101101011: color_data = 12'b111100001111;
20'b01101100010101101100: color_data = 12'b111100001111;
20'b01101100010101101101: color_data = 12'b111100001111;
20'b01101100010101101110: color_data = 12'b111100001111;
20'b01101100010101101111: color_data = 12'b111100001111;
20'b01101100010101110000: color_data = 12'b111100001111;
20'b01101100010101110001: color_data = 12'b111100001111;
20'b01101100010101110010: color_data = 12'b111100001111;
20'b01101100010101110011: color_data = 12'b111100001111;
20'b01101100010101110100: color_data = 12'b111100001111;
20'b01101100010101111000: color_data = 12'b111100000000;
20'b01101100010101111001: color_data = 12'b111100000000;
20'b01101100010101111010: color_data = 12'b111100000000;
20'b01101100010101111011: color_data = 12'b111100000000;
20'b01101100010101111100: color_data = 12'b111100000000;
20'b01101100010101111101: color_data = 12'b111100000000;
20'b01101100010101111110: color_data = 12'b111100000000;
20'b01101100010101111111: color_data = 12'b111100000000;
20'b01101100010110000000: color_data = 12'b111100000000;
20'b01101100010110000001: color_data = 12'b111100000000;
20'b01101100010110000010: color_data = 12'b111100000000;
20'b01101100010110000011: color_data = 12'b111100000000;
20'b01101100010110000100: color_data = 12'b111100000000;
20'b01101100010110000101: color_data = 12'b111100000000;
20'b01101100010110000110: color_data = 12'b111100000000;
20'b01101100010110000111: color_data = 12'b111100000000;
20'b01101100010110001000: color_data = 12'b111100000000;
20'b01101100010110001001: color_data = 12'b111100000000;
20'b01101100010110001101: color_data = 12'b111100000000;
20'b01101100010110001110: color_data = 12'b111100000000;
20'b01101100010110001111: color_data = 12'b111100000000;
20'b01101100010110010000: color_data = 12'b111100000000;
20'b01101100010110010001: color_data = 12'b111100000000;
20'b01101100010110010010: color_data = 12'b111100000000;
20'b01101100010110010011: color_data = 12'b111100000000;
20'b01101100010110010100: color_data = 12'b111100000000;
20'b01101100010110010101: color_data = 12'b111100000000;
20'b01101100010110010110: color_data = 12'b111100000000;
20'b01101100010110010111: color_data = 12'b111100000000;
20'b01101100010110011000: color_data = 12'b111100000000;
20'b01101100010110011001: color_data = 12'b111100000000;
20'b01101100010110011010: color_data = 12'b111100000000;
20'b01101100010110011011: color_data = 12'b111100000000;
20'b01101100010110011100: color_data = 12'b111100000000;
20'b01101100010110011101: color_data = 12'b111100000000;
20'b01101100010110011110: color_data = 12'b111100000000;
20'b01101100100011111010: color_data = 12'b111101110000;
20'b01101100100011111011: color_data = 12'b111101110000;
20'b01101100100011111100: color_data = 12'b111101110000;
20'b01101100100011111101: color_data = 12'b111101110000;
20'b01101100100011111110: color_data = 12'b111101110000;
20'b01101100100011111111: color_data = 12'b111101110000;
20'b01101100100100000000: color_data = 12'b111101110000;
20'b01101100100100000001: color_data = 12'b111101110000;
20'b01101100100100000010: color_data = 12'b111101110000;
20'b01101100100100000011: color_data = 12'b111101110000;
20'b01101100100100000100: color_data = 12'b111101110000;
20'b01101100100100000101: color_data = 12'b111101110000;
20'b01101100100100000110: color_data = 12'b111101110000;
20'b01101100100100000111: color_data = 12'b111101110000;
20'b01101100100100001000: color_data = 12'b111101110000;
20'b01101100100100001001: color_data = 12'b111101110000;
20'b01101100100100001010: color_data = 12'b111101110000;
20'b01101100100100001011: color_data = 12'b111101110000;
20'b01101100100100001111: color_data = 12'b111101110000;
20'b01101100100100010000: color_data = 12'b111101110000;
20'b01101100100100010001: color_data = 12'b111101110000;
20'b01101100100100010010: color_data = 12'b111101110000;
20'b01101100100100010011: color_data = 12'b111101110000;
20'b01101100100100010100: color_data = 12'b111101110000;
20'b01101100100100010101: color_data = 12'b111101110000;
20'b01101100100100010110: color_data = 12'b111101110000;
20'b01101100100100010111: color_data = 12'b111101110000;
20'b01101100100100011000: color_data = 12'b111101110000;
20'b01101100100100011001: color_data = 12'b111101110000;
20'b01101100100100011010: color_data = 12'b111101110000;
20'b01101100100100011011: color_data = 12'b111101110000;
20'b01101100100100011100: color_data = 12'b111101110000;
20'b01101100100100011101: color_data = 12'b111101110000;
20'b01101100100100011110: color_data = 12'b111101110000;
20'b01101100100100011111: color_data = 12'b111101110000;
20'b01101100100100100000: color_data = 12'b111101110000;
20'b01101100100100100100: color_data = 12'b111101110000;
20'b01101100100100100101: color_data = 12'b111101110000;
20'b01101100100100100110: color_data = 12'b111101110000;
20'b01101100100100100111: color_data = 12'b111101110000;
20'b01101100100100101000: color_data = 12'b111101110000;
20'b01101100100100101001: color_data = 12'b111101110000;
20'b01101100100100101010: color_data = 12'b111101110000;
20'b01101100100100101011: color_data = 12'b111101110000;
20'b01101100100100101100: color_data = 12'b111101110000;
20'b01101100100100101101: color_data = 12'b111101110000;
20'b01101100100100101110: color_data = 12'b111101110000;
20'b01101100100100101111: color_data = 12'b111101110000;
20'b01101100100100110000: color_data = 12'b111101110000;
20'b01101100100100110001: color_data = 12'b111101110000;
20'b01101100100100110010: color_data = 12'b111101110000;
20'b01101100100100110011: color_data = 12'b111101110000;
20'b01101100100100110100: color_data = 12'b111101110000;
20'b01101100100100110101: color_data = 12'b111101110000;
20'b01101100100100111001: color_data = 12'b111101110000;
20'b01101100100100111010: color_data = 12'b111101110000;
20'b01101100100100111011: color_data = 12'b111101110000;
20'b01101100100100111100: color_data = 12'b111101110000;
20'b01101100100100111101: color_data = 12'b111101110000;
20'b01101100100100111110: color_data = 12'b111101110000;
20'b01101100100100111111: color_data = 12'b111101110000;
20'b01101100100101000000: color_data = 12'b111101110000;
20'b01101100100101000001: color_data = 12'b111101110000;
20'b01101100100101000010: color_data = 12'b111101110000;
20'b01101100100101000011: color_data = 12'b111101110000;
20'b01101100100101000100: color_data = 12'b111101110000;
20'b01101100100101000101: color_data = 12'b111101110000;
20'b01101100100101000110: color_data = 12'b111101110000;
20'b01101100100101000111: color_data = 12'b111101110000;
20'b01101100100101001000: color_data = 12'b111101110000;
20'b01101100100101001001: color_data = 12'b111101110000;
20'b01101100100101001010: color_data = 12'b111101110000;
20'b01101100100101001110: color_data = 12'b000011110000;
20'b01101100100101001111: color_data = 12'b000011110000;
20'b01101100100101010000: color_data = 12'b000011110000;
20'b01101100100101010001: color_data = 12'b000011110000;
20'b01101100100101010010: color_data = 12'b000011110000;
20'b01101100100101010011: color_data = 12'b000011110000;
20'b01101100100101010100: color_data = 12'b000011110000;
20'b01101100100101010101: color_data = 12'b000011110000;
20'b01101100100101010110: color_data = 12'b000011110000;
20'b01101100100101010111: color_data = 12'b000011110000;
20'b01101100100101011000: color_data = 12'b000011110000;
20'b01101100100101011001: color_data = 12'b000011110000;
20'b01101100100101011010: color_data = 12'b000011110000;
20'b01101100100101011011: color_data = 12'b000011110000;
20'b01101100100101011100: color_data = 12'b000011110000;
20'b01101100100101011101: color_data = 12'b000011110000;
20'b01101100100101011110: color_data = 12'b000011110000;
20'b01101100100101011111: color_data = 12'b000011110000;
20'b01101100100101100011: color_data = 12'b111100001111;
20'b01101100100101100100: color_data = 12'b111100001111;
20'b01101100100101100101: color_data = 12'b111100001111;
20'b01101100100101100110: color_data = 12'b111100001111;
20'b01101100100101100111: color_data = 12'b111100001111;
20'b01101100100101101000: color_data = 12'b111100001111;
20'b01101100100101101001: color_data = 12'b111100001111;
20'b01101100100101101010: color_data = 12'b111100001111;
20'b01101100100101101011: color_data = 12'b111100001111;
20'b01101100100101101100: color_data = 12'b111100001111;
20'b01101100100101101101: color_data = 12'b111100001111;
20'b01101100100101101110: color_data = 12'b111100001111;
20'b01101100100101101111: color_data = 12'b111100001111;
20'b01101100100101110000: color_data = 12'b111100001111;
20'b01101100100101110001: color_data = 12'b111100001111;
20'b01101100100101110010: color_data = 12'b111100001111;
20'b01101100100101110011: color_data = 12'b111100001111;
20'b01101100100101110100: color_data = 12'b111100001111;
20'b01101100100101111000: color_data = 12'b111100000000;
20'b01101100100101111001: color_data = 12'b111100000000;
20'b01101100100101111010: color_data = 12'b111100000000;
20'b01101100100101111011: color_data = 12'b111100000000;
20'b01101100100101111100: color_data = 12'b111100000000;
20'b01101100100101111101: color_data = 12'b111100000000;
20'b01101100100101111110: color_data = 12'b111100000000;
20'b01101100100101111111: color_data = 12'b111100000000;
20'b01101100100110000000: color_data = 12'b111100000000;
20'b01101100100110000001: color_data = 12'b111100000000;
20'b01101100100110000010: color_data = 12'b111100000000;
20'b01101100100110000011: color_data = 12'b111100000000;
20'b01101100100110000100: color_data = 12'b111100000000;
20'b01101100100110000101: color_data = 12'b111100000000;
20'b01101100100110000110: color_data = 12'b111100000000;
20'b01101100100110000111: color_data = 12'b111100000000;
20'b01101100100110001000: color_data = 12'b111100000000;
20'b01101100100110001001: color_data = 12'b111100000000;
20'b01101100100110001101: color_data = 12'b111100000000;
20'b01101100100110001110: color_data = 12'b111100000000;
20'b01101100100110001111: color_data = 12'b111100000000;
20'b01101100100110010000: color_data = 12'b111100000000;
20'b01101100100110010001: color_data = 12'b111100000000;
20'b01101100100110010010: color_data = 12'b111100000000;
20'b01101100100110010011: color_data = 12'b111100000000;
20'b01101100100110010100: color_data = 12'b111100000000;
20'b01101100100110010101: color_data = 12'b111100000000;
20'b01101100100110010110: color_data = 12'b111100000000;
20'b01101100100110010111: color_data = 12'b111100000000;
20'b01101100100110011000: color_data = 12'b111100000000;
20'b01101100100110011001: color_data = 12'b111100000000;
20'b01101100100110011010: color_data = 12'b111100000000;
20'b01101100100110011011: color_data = 12'b111100000000;
20'b01101100100110011100: color_data = 12'b111100000000;
20'b01101100100110011101: color_data = 12'b111100000000;
20'b01101100100110011110: color_data = 12'b111100000000;
20'b01101100110011111010: color_data = 12'b111101110000;
20'b01101100110011111011: color_data = 12'b111101110000;
20'b01101100110011111100: color_data = 12'b111101110000;
20'b01101100110011111101: color_data = 12'b111101110000;
20'b01101100110011111110: color_data = 12'b111101110000;
20'b01101100110011111111: color_data = 12'b111101110000;
20'b01101100110100000000: color_data = 12'b111101110000;
20'b01101100110100000001: color_data = 12'b111101110000;
20'b01101100110100000010: color_data = 12'b111101110000;
20'b01101100110100000011: color_data = 12'b111101110000;
20'b01101100110100000100: color_data = 12'b111101110000;
20'b01101100110100000101: color_data = 12'b111101110000;
20'b01101100110100000110: color_data = 12'b111101110000;
20'b01101100110100000111: color_data = 12'b111101110000;
20'b01101100110100001000: color_data = 12'b111101110000;
20'b01101100110100001001: color_data = 12'b111101110000;
20'b01101100110100001010: color_data = 12'b111101110000;
20'b01101100110100001011: color_data = 12'b111101110000;
20'b01101100110100001111: color_data = 12'b111101110000;
20'b01101100110100010000: color_data = 12'b111101110000;
20'b01101100110100010001: color_data = 12'b111101110000;
20'b01101100110100010010: color_data = 12'b111101110000;
20'b01101100110100010011: color_data = 12'b111101110000;
20'b01101100110100010100: color_data = 12'b111101110000;
20'b01101100110100010101: color_data = 12'b111101110000;
20'b01101100110100010110: color_data = 12'b111101110000;
20'b01101100110100010111: color_data = 12'b111101110000;
20'b01101100110100011000: color_data = 12'b111101110000;
20'b01101100110100011001: color_data = 12'b111101110000;
20'b01101100110100011010: color_data = 12'b111101110000;
20'b01101100110100011011: color_data = 12'b111101110000;
20'b01101100110100011100: color_data = 12'b111101110000;
20'b01101100110100011101: color_data = 12'b111101110000;
20'b01101100110100011110: color_data = 12'b111101110000;
20'b01101100110100011111: color_data = 12'b111101110000;
20'b01101100110100100000: color_data = 12'b111101110000;
20'b01101100110100100100: color_data = 12'b111101110000;
20'b01101100110100100101: color_data = 12'b111101110000;
20'b01101100110100100110: color_data = 12'b111101110000;
20'b01101100110100100111: color_data = 12'b111101110000;
20'b01101100110100101000: color_data = 12'b111101110000;
20'b01101100110100101001: color_data = 12'b111101110000;
20'b01101100110100101010: color_data = 12'b111101110000;
20'b01101100110100101011: color_data = 12'b111101110000;
20'b01101100110100101100: color_data = 12'b111101110000;
20'b01101100110100101101: color_data = 12'b111101110000;
20'b01101100110100101110: color_data = 12'b111101110000;
20'b01101100110100101111: color_data = 12'b111101110000;
20'b01101100110100110000: color_data = 12'b111101110000;
20'b01101100110100110001: color_data = 12'b111101110000;
20'b01101100110100110010: color_data = 12'b111101110000;
20'b01101100110100110011: color_data = 12'b111101110000;
20'b01101100110100110100: color_data = 12'b111101110000;
20'b01101100110100110101: color_data = 12'b111101110000;
20'b01101100110100111001: color_data = 12'b111101110000;
20'b01101100110100111010: color_data = 12'b111101110000;
20'b01101100110100111011: color_data = 12'b111101110000;
20'b01101100110100111100: color_data = 12'b111101110000;
20'b01101100110100111101: color_data = 12'b111101110000;
20'b01101100110100111110: color_data = 12'b111101110000;
20'b01101100110100111111: color_data = 12'b111101110000;
20'b01101100110101000000: color_data = 12'b111101110000;
20'b01101100110101000001: color_data = 12'b111101110000;
20'b01101100110101000010: color_data = 12'b111101110000;
20'b01101100110101000011: color_data = 12'b111101110000;
20'b01101100110101000100: color_data = 12'b111101110000;
20'b01101100110101000101: color_data = 12'b111101110000;
20'b01101100110101000110: color_data = 12'b111101110000;
20'b01101100110101000111: color_data = 12'b111101110000;
20'b01101100110101001000: color_data = 12'b111101110000;
20'b01101100110101001001: color_data = 12'b111101110000;
20'b01101100110101001010: color_data = 12'b111101110000;
20'b01101100110101001110: color_data = 12'b000011110000;
20'b01101100110101001111: color_data = 12'b000011110000;
20'b01101100110101010000: color_data = 12'b000011110000;
20'b01101100110101010001: color_data = 12'b000011110000;
20'b01101100110101010010: color_data = 12'b000011110000;
20'b01101100110101010011: color_data = 12'b000011110000;
20'b01101100110101010100: color_data = 12'b000011110000;
20'b01101100110101010101: color_data = 12'b000011110000;
20'b01101100110101010110: color_data = 12'b000011110000;
20'b01101100110101010111: color_data = 12'b000011110000;
20'b01101100110101011000: color_data = 12'b000011110000;
20'b01101100110101011001: color_data = 12'b000011110000;
20'b01101100110101011010: color_data = 12'b000011110000;
20'b01101100110101011011: color_data = 12'b000011110000;
20'b01101100110101011100: color_data = 12'b000011110000;
20'b01101100110101011101: color_data = 12'b000011110000;
20'b01101100110101011110: color_data = 12'b000011110000;
20'b01101100110101011111: color_data = 12'b000011110000;
20'b01101100110101100011: color_data = 12'b111100001111;
20'b01101100110101100100: color_data = 12'b111100001111;
20'b01101100110101100101: color_data = 12'b111100001111;
20'b01101100110101100110: color_data = 12'b111100001111;
20'b01101100110101100111: color_data = 12'b111100001111;
20'b01101100110101101000: color_data = 12'b111100001111;
20'b01101100110101101001: color_data = 12'b111100001111;
20'b01101100110101101010: color_data = 12'b111100001111;
20'b01101100110101101011: color_data = 12'b111100001111;
20'b01101100110101101100: color_data = 12'b111100001111;
20'b01101100110101101101: color_data = 12'b111100001111;
20'b01101100110101101110: color_data = 12'b111100001111;
20'b01101100110101101111: color_data = 12'b111100001111;
20'b01101100110101110000: color_data = 12'b111100001111;
20'b01101100110101110001: color_data = 12'b111100001111;
20'b01101100110101110010: color_data = 12'b111100001111;
20'b01101100110101110011: color_data = 12'b111100001111;
20'b01101100110101110100: color_data = 12'b111100001111;
20'b01101100110101111000: color_data = 12'b111100000000;
20'b01101100110101111001: color_data = 12'b111100000000;
20'b01101100110101111010: color_data = 12'b111100000000;
20'b01101100110101111011: color_data = 12'b111100000000;
20'b01101100110101111100: color_data = 12'b111100000000;
20'b01101100110101111101: color_data = 12'b111100000000;
20'b01101100110101111110: color_data = 12'b111100000000;
20'b01101100110101111111: color_data = 12'b111100000000;
20'b01101100110110000000: color_data = 12'b111100000000;
20'b01101100110110000001: color_data = 12'b111100000000;
20'b01101100110110000010: color_data = 12'b111100000000;
20'b01101100110110000011: color_data = 12'b111100000000;
20'b01101100110110000100: color_data = 12'b111100000000;
20'b01101100110110000101: color_data = 12'b111100000000;
20'b01101100110110000110: color_data = 12'b111100000000;
20'b01101100110110000111: color_data = 12'b111100000000;
20'b01101100110110001000: color_data = 12'b111100000000;
20'b01101100110110001001: color_data = 12'b111100000000;
20'b01101100110110001101: color_data = 12'b111100000000;
20'b01101100110110001110: color_data = 12'b111100000000;
20'b01101100110110001111: color_data = 12'b111100000000;
20'b01101100110110010000: color_data = 12'b111100000000;
20'b01101100110110010001: color_data = 12'b111100000000;
20'b01101100110110010010: color_data = 12'b111100000000;
20'b01101100110110010011: color_data = 12'b111100000000;
20'b01101100110110010100: color_data = 12'b111100000000;
20'b01101100110110010101: color_data = 12'b111100000000;
20'b01101100110110010110: color_data = 12'b111100000000;
20'b01101100110110010111: color_data = 12'b111100000000;
20'b01101100110110011000: color_data = 12'b111100000000;
20'b01101100110110011001: color_data = 12'b111100000000;
20'b01101100110110011010: color_data = 12'b111100000000;
20'b01101100110110011011: color_data = 12'b111100000000;
20'b01101100110110011100: color_data = 12'b111100000000;
20'b01101100110110011101: color_data = 12'b111100000000;
20'b01101100110110011110: color_data = 12'b111100000000;
20'b01101101000011111010: color_data = 12'b111101110000;
20'b01101101000011111011: color_data = 12'b111101110000;
20'b01101101000011111100: color_data = 12'b111101110000;
20'b01101101000011111101: color_data = 12'b111101110000;
20'b01101101000011111110: color_data = 12'b111101110000;
20'b01101101000011111111: color_data = 12'b111101110000;
20'b01101101000100000000: color_data = 12'b111101110000;
20'b01101101000100000001: color_data = 12'b111101110000;
20'b01101101000100000010: color_data = 12'b111101110000;
20'b01101101000100000011: color_data = 12'b111101110000;
20'b01101101000100000100: color_data = 12'b111101110000;
20'b01101101000100000101: color_data = 12'b111101110000;
20'b01101101000100000110: color_data = 12'b111101110000;
20'b01101101000100000111: color_data = 12'b111101110000;
20'b01101101000100001000: color_data = 12'b111101110000;
20'b01101101000100001001: color_data = 12'b111101110000;
20'b01101101000100001010: color_data = 12'b111101110000;
20'b01101101000100001011: color_data = 12'b111101110000;
20'b01101101000100001111: color_data = 12'b111101110000;
20'b01101101000100010000: color_data = 12'b111101110000;
20'b01101101000100010001: color_data = 12'b111101110000;
20'b01101101000100010010: color_data = 12'b111101110000;
20'b01101101000100010011: color_data = 12'b111101110000;
20'b01101101000100010100: color_data = 12'b111101110000;
20'b01101101000100010101: color_data = 12'b111101110000;
20'b01101101000100010110: color_data = 12'b111101110000;
20'b01101101000100010111: color_data = 12'b111101110000;
20'b01101101000100011000: color_data = 12'b111101110000;
20'b01101101000100011001: color_data = 12'b111101110000;
20'b01101101000100011010: color_data = 12'b111101110000;
20'b01101101000100011011: color_data = 12'b111101110000;
20'b01101101000100011100: color_data = 12'b111101110000;
20'b01101101000100011101: color_data = 12'b111101110000;
20'b01101101000100011110: color_data = 12'b111101110000;
20'b01101101000100011111: color_data = 12'b111101110000;
20'b01101101000100100000: color_data = 12'b111101110000;
20'b01101101000100100100: color_data = 12'b111101110000;
20'b01101101000100100101: color_data = 12'b111101110000;
20'b01101101000100100110: color_data = 12'b111101110000;
20'b01101101000100100111: color_data = 12'b111101110000;
20'b01101101000100101000: color_data = 12'b111101110000;
20'b01101101000100101001: color_data = 12'b111101110000;
20'b01101101000100101010: color_data = 12'b111101110000;
20'b01101101000100101011: color_data = 12'b111101110000;
20'b01101101000100101100: color_data = 12'b111101110000;
20'b01101101000100101101: color_data = 12'b111101110000;
20'b01101101000100101110: color_data = 12'b111101110000;
20'b01101101000100101111: color_data = 12'b111101110000;
20'b01101101000100110000: color_data = 12'b111101110000;
20'b01101101000100110001: color_data = 12'b111101110000;
20'b01101101000100110010: color_data = 12'b111101110000;
20'b01101101000100110011: color_data = 12'b111101110000;
20'b01101101000100110100: color_data = 12'b111101110000;
20'b01101101000100110101: color_data = 12'b111101110000;
20'b01101101000100111001: color_data = 12'b111101110000;
20'b01101101000100111010: color_data = 12'b111101110000;
20'b01101101000100111011: color_data = 12'b111101110000;
20'b01101101000100111100: color_data = 12'b111101110000;
20'b01101101000100111101: color_data = 12'b111101110000;
20'b01101101000100111110: color_data = 12'b111101110000;
20'b01101101000100111111: color_data = 12'b111101110000;
20'b01101101000101000000: color_data = 12'b111101110000;
20'b01101101000101000001: color_data = 12'b111101110000;
20'b01101101000101000010: color_data = 12'b111101110000;
20'b01101101000101000011: color_data = 12'b111101110000;
20'b01101101000101000100: color_data = 12'b111101110000;
20'b01101101000101000101: color_data = 12'b111101110000;
20'b01101101000101000110: color_data = 12'b111101110000;
20'b01101101000101000111: color_data = 12'b111101110000;
20'b01101101000101001000: color_data = 12'b111101110000;
20'b01101101000101001001: color_data = 12'b111101110000;
20'b01101101000101001010: color_data = 12'b111101110000;
20'b01101101000101001110: color_data = 12'b000011110000;
20'b01101101000101001111: color_data = 12'b000011110000;
20'b01101101000101010000: color_data = 12'b000011110000;
20'b01101101000101010001: color_data = 12'b000011110000;
20'b01101101000101010010: color_data = 12'b000011110000;
20'b01101101000101010011: color_data = 12'b000011110000;
20'b01101101000101010100: color_data = 12'b000011110000;
20'b01101101000101010101: color_data = 12'b000011110000;
20'b01101101000101010110: color_data = 12'b000011110000;
20'b01101101000101010111: color_data = 12'b000011110000;
20'b01101101000101011000: color_data = 12'b000011110000;
20'b01101101000101011001: color_data = 12'b000011110000;
20'b01101101000101011010: color_data = 12'b000011110000;
20'b01101101000101011011: color_data = 12'b000011110000;
20'b01101101000101011100: color_data = 12'b000011110000;
20'b01101101000101011101: color_data = 12'b000011110000;
20'b01101101000101011110: color_data = 12'b000011110000;
20'b01101101000101011111: color_data = 12'b000011110000;
20'b01101101000101100011: color_data = 12'b111100001111;
20'b01101101000101100100: color_data = 12'b111100001111;
20'b01101101000101100101: color_data = 12'b111100001111;
20'b01101101000101100110: color_data = 12'b111100001111;
20'b01101101000101100111: color_data = 12'b111100001111;
20'b01101101000101101000: color_data = 12'b111100001111;
20'b01101101000101101001: color_data = 12'b111100001111;
20'b01101101000101101010: color_data = 12'b111100001111;
20'b01101101000101101011: color_data = 12'b111100001111;
20'b01101101000101101100: color_data = 12'b111100001111;
20'b01101101000101101101: color_data = 12'b111100001111;
20'b01101101000101101110: color_data = 12'b111100001111;
20'b01101101000101101111: color_data = 12'b111100001111;
20'b01101101000101110000: color_data = 12'b111100001111;
20'b01101101000101110001: color_data = 12'b111100001111;
20'b01101101000101110010: color_data = 12'b111100001111;
20'b01101101000101110011: color_data = 12'b111100001111;
20'b01101101000101110100: color_data = 12'b111100001111;
20'b01101101000101111000: color_data = 12'b111100000000;
20'b01101101000101111001: color_data = 12'b111100000000;
20'b01101101000101111010: color_data = 12'b111100000000;
20'b01101101000101111011: color_data = 12'b111100000000;
20'b01101101000101111100: color_data = 12'b111100000000;
20'b01101101000101111101: color_data = 12'b111100000000;
20'b01101101000101111110: color_data = 12'b111100000000;
20'b01101101000101111111: color_data = 12'b111100000000;
20'b01101101000110000000: color_data = 12'b111100000000;
20'b01101101000110000001: color_data = 12'b111100000000;
20'b01101101000110000010: color_data = 12'b111100000000;
20'b01101101000110000011: color_data = 12'b111100000000;
20'b01101101000110000100: color_data = 12'b111100000000;
20'b01101101000110000101: color_data = 12'b111100000000;
20'b01101101000110000110: color_data = 12'b111100000000;
20'b01101101000110000111: color_data = 12'b111100000000;
20'b01101101000110001000: color_data = 12'b111100000000;
20'b01101101000110001001: color_data = 12'b111100000000;
20'b01101101000110001101: color_data = 12'b111100000000;
20'b01101101000110001110: color_data = 12'b111100000000;
20'b01101101000110001111: color_data = 12'b111100000000;
20'b01101101000110010000: color_data = 12'b111100000000;
20'b01101101000110010001: color_data = 12'b111100000000;
20'b01101101000110010010: color_data = 12'b111100000000;
20'b01101101000110010011: color_data = 12'b111100000000;
20'b01101101000110010100: color_data = 12'b111100000000;
20'b01101101000110010101: color_data = 12'b111100000000;
20'b01101101000110010110: color_data = 12'b111100000000;
20'b01101101000110010111: color_data = 12'b111100000000;
20'b01101101000110011000: color_data = 12'b111100000000;
20'b01101101000110011001: color_data = 12'b111100000000;
20'b01101101000110011010: color_data = 12'b111100000000;
20'b01101101000110011011: color_data = 12'b111100000000;
20'b01101101000110011100: color_data = 12'b111100000000;
20'b01101101000110011101: color_data = 12'b111100000000;
20'b01101101000110011110: color_data = 12'b111100000000;
20'b01101101010011111010: color_data = 12'b111101110000;
20'b01101101010011111011: color_data = 12'b111101110000;
20'b01101101010011111100: color_data = 12'b111101110000;
20'b01101101010011111101: color_data = 12'b111101110000;
20'b01101101010011111110: color_data = 12'b111101110000;
20'b01101101010011111111: color_data = 12'b111101110000;
20'b01101101010100000000: color_data = 12'b111101110000;
20'b01101101010100000001: color_data = 12'b111101110000;
20'b01101101010100000010: color_data = 12'b111101110000;
20'b01101101010100000011: color_data = 12'b111101110000;
20'b01101101010100000100: color_data = 12'b111101110000;
20'b01101101010100000101: color_data = 12'b111101110000;
20'b01101101010100000110: color_data = 12'b111101110000;
20'b01101101010100000111: color_data = 12'b111101110000;
20'b01101101010100001000: color_data = 12'b111101110000;
20'b01101101010100001001: color_data = 12'b111101110000;
20'b01101101010100001010: color_data = 12'b111101110000;
20'b01101101010100001011: color_data = 12'b111101110000;
20'b01101101010100001111: color_data = 12'b111101110000;
20'b01101101010100010000: color_data = 12'b111101110000;
20'b01101101010100010001: color_data = 12'b111101110000;
20'b01101101010100010010: color_data = 12'b111101110000;
20'b01101101010100010011: color_data = 12'b111101110000;
20'b01101101010100010100: color_data = 12'b111101110000;
20'b01101101010100010101: color_data = 12'b111101110000;
20'b01101101010100010110: color_data = 12'b111101110000;
20'b01101101010100010111: color_data = 12'b111101110000;
20'b01101101010100011000: color_data = 12'b111101110000;
20'b01101101010100011001: color_data = 12'b111101110000;
20'b01101101010100011010: color_data = 12'b111101110000;
20'b01101101010100011011: color_data = 12'b111101110000;
20'b01101101010100011100: color_data = 12'b111101110000;
20'b01101101010100011101: color_data = 12'b111101110000;
20'b01101101010100011110: color_data = 12'b111101110000;
20'b01101101010100011111: color_data = 12'b111101110000;
20'b01101101010100100000: color_data = 12'b111101110000;
20'b01101101010100100100: color_data = 12'b111101110000;
20'b01101101010100100101: color_data = 12'b111101110000;
20'b01101101010100100110: color_data = 12'b111101110000;
20'b01101101010100100111: color_data = 12'b111101110000;
20'b01101101010100101000: color_data = 12'b111101110000;
20'b01101101010100101001: color_data = 12'b111101110000;
20'b01101101010100101010: color_data = 12'b111101110000;
20'b01101101010100101011: color_data = 12'b111101110000;
20'b01101101010100101100: color_data = 12'b111101110000;
20'b01101101010100101101: color_data = 12'b111101110000;
20'b01101101010100101110: color_data = 12'b111101110000;
20'b01101101010100101111: color_data = 12'b111101110000;
20'b01101101010100110000: color_data = 12'b111101110000;
20'b01101101010100110001: color_data = 12'b111101110000;
20'b01101101010100110010: color_data = 12'b111101110000;
20'b01101101010100110011: color_data = 12'b111101110000;
20'b01101101010100110100: color_data = 12'b111101110000;
20'b01101101010100110101: color_data = 12'b111101110000;
20'b01101101010100111001: color_data = 12'b111101110000;
20'b01101101010100111010: color_data = 12'b111101110000;
20'b01101101010100111011: color_data = 12'b111101110000;
20'b01101101010100111100: color_data = 12'b111101110000;
20'b01101101010100111101: color_data = 12'b111101110000;
20'b01101101010100111110: color_data = 12'b111101110000;
20'b01101101010100111111: color_data = 12'b111101110000;
20'b01101101010101000000: color_data = 12'b111101110000;
20'b01101101010101000001: color_data = 12'b111101110000;
20'b01101101010101000010: color_data = 12'b111101110000;
20'b01101101010101000011: color_data = 12'b111101110000;
20'b01101101010101000100: color_data = 12'b111101110000;
20'b01101101010101000101: color_data = 12'b111101110000;
20'b01101101010101000110: color_data = 12'b111101110000;
20'b01101101010101000111: color_data = 12'b111101110000;
20'b01101101010101001000: color_data = 12'b111101110000;
20'b01101101010101001001: color_data = 12'b111101110000;
20'b01101101010101001010: color_data = 12'b111101110000;
20'b01101101010101001110: color_data = 12'b000011110000;
20'b01101101010101001111: color_data = 12'b000011110000;
20'b01101101010101010000: color_data = 12'b000011110000;
20'b01101101010101010001: color_data = 12'b000011110000;
20'b01101101010101010010: color_data = 12'b000011110000;
20'b01101101010101010011: color_data = 12'b000011110000;
20'b01101101010101010100: color_data = 12'b000011110000;
20'b01101101010101010101: color_data = 12'b000011110000;
20'b01101101010101010110: color_data = 12'b000011110000;
20'b01101101010101010111: color_data = 12'b000011110000;
20'b01101101010101011000: color_data = 12'b000011110000;
20'b01101101010101011001: color_data = 12'b000011110000;
20'b01101101010101011010: color_data = 12'b000011110000;
20'b01101101010101011011: color_data = 12'b000011110000;
20'b01101101010101011100: color_data = 12'b000011110000;
20'b01101101010101011101: color_data = 12'b000011110000;
20'b01101101010101011110: color_data = 12'b000011110000;
20'b01101101010101011111: color_data = 12'b000011110000;
20'b01101101010101100011: color_data = 12'b111100001111;
20'b01101101010101100100: color_data = 12'b111100001111;
20'b01101101010101100101: color_data = 12'b111100001111;
20'b01101101010101100110: color_data = 12'b111100001111;
20'b01101101010101100111: color_data = 12'b111100001111;
20'b01101101010101101000: color_data = 12'b111100001111;
20'b01101101010101101001: color_data = 12'b111100001111;
20'b01101101010101101010: color_data = 12'b111100001111;
20'b01101101010101101011: color_data = 12'b111100001111;
20'b01101101010101101100: color_data = 12'b111100001111;
20'b01101101010101101101: color_data = 12'b111100001111;
20'b01101101010101101110: color_data = 12'b111100001111;
20'b01101101010101101111: color_data = 12'b111100001111;
20'b01101101010101110000: color_data = 12'b111100001111;
20'b01101101010101110001: color_data = 12'b111100001111;
20'b01101101010101110010: color_data = 12'b111100001111;
20'b01101101010101110011: color_data = 12'b111100001111;
20'b01101101010101110100: color_data = 12'b111100001111;
20'b01101101010101111000: color_data = 12'b111100000000;
20'b01101101010101111001: color_data = 12'b111100000000;
20'b01101101010101111010: color_data = 12'b111100000000;
20'b01101101010101111011: color_data = 12'b111100000000;
20'b01101101010101111100: color_data = 12'b111100000000;
20'b01101101010101111101: color_data = 12'b111100000000;
20'b01101101010101111110: color_data = 12'b111100000000;
20'b01101101010101111111: color_data = 12'b111100000000;
20'b01101101010110000000: color_data = 12'b111100000000;
20'b01101101010110000001: color_data = 12'b111100000000;
20'b01101101010110000010: color_data = 12'b111100000000;
20'b01101101010110000011: color_data = 12'b111100000000;
20'b01101101010110000100: color_data = 12'b111100000000;
20'b01101101010110000101: color_data = 12'b111100000000;
20'b01101101010110000110: color_data = 12'b111100000000;
20'b01101101010110000111: color_data = 12'b111100000000;
20'b01101101010110001000: color_data = 12'b111100000000;
20'b01101101010110001001: color_data = 12'b111100000000;
20'b01101101010110001101: color_data = 12'b111100000000;
20'b01101101010110001110: color_data = 12'b111100000000;
20'b01101101010110001111: color_data = 12'b111100000000;
20'b01101101010110010000: color_data = 12'b111100000000;
20'b01101101010110010001: color_data = 12'b111100000000;
20'b01101101010110010010: color_data = 12'b111100000000;
20'b01101101010110010011: color_data = 12'b111100000000;
20'b01101101010110010100: color_data = 12'b111100000000;
20'b01101101010110010101: color_data = 12'b111100000000;
20'b01101101010110010110: color_data = 12'b111100000000;
20'b01101101010110010111: color_data = 12'b111100000000;
20'b01101101010110011000: color_data = 12'b111100000000;
20'b01101101010110011001: color_data = 12'b111100000000;
20'b01101101010110011010: color_data = 12'b111100000000;
20'b01101101010110011011: color_data = 12'b111100000000;
20'b01101101010110011100: color_data = 12'b111100000000;
20'b01101101010110011101: color_data = 12'b111100000000;
20'b01101101010110011110: color_data = 12'b111100000000;
20'b01101101100011111010: color_data = 12'b111101110000;
20'b01101101100011111011: color_data = 12'b111101110000;
20'b01101101100011111100: color_data = 12'b111101110000;
20'b01101101100011111101: color_data = 12'b111101110000;
20'b01101101100011111110: color_data = 12'b111101110000;
20'b01101101100011111111: color_data = 12'b111101110000;
20'b01101101100100000000: color_data = 12'b111101110000;
20'b01101101100100000001: color_data = 12'b111101110000;
20'b01101101100100000010: color_data = 12'b111101110000;
20'b01101101100100000011: color_data = 12'b111101110000;
20'b01101101100100000100: color_data = 12'b111101110000;
20'b01101101100100000101: color_data = 12'b111101110000;
20'b01101101100100000110: color_data = 12'b111101110000;
20'b01101101100100000111: color_data = 12'b111101110000;
20'b01101101100100001000: color_data = 12'b111101110000;
20'b01101101100100001001: color_data = 12'b111101110000;
20'b01101101100100001010: color_data = 12'b111101110000;
20'b01101101100100001011: color_data = 12'b111101110000;
20'b01101101100100001111: color_data = 12'b111101110000;
20'b01101101100100010000: color_data = 12'b111101110000;
20'b01101101100100010001: color_data = 12'b111101110000;
20'b01101101100100010010: color_data = 12'b111101110000;
20'b01101101100100010011: color_data = 12'b111101110000;
20'b01101101100100010100: color_data = 12'b111101110000;
20'b01101101100100010101: color_data = 12'b111101110000;
20'b01101101100100010110: color_data = 12'b111101110000;
20'b01101101100100010111: color_data = 12'b111101110000;
20'b01101101100100011000: color_data = 12'b111101110000;
20'b01101101100100011001: color_data = 12'b111101110000;
20'b01101101100100011010: color_data = 12'b111101110000;
20'b01101101100100011011: color_data = 12'b111101110000;
20'b01101101100100011100: color_data = 12'b111101110000;
20'b01101101100100011101: color_data = 12'b111101110000;
20'b01101101100100011110: color_data = 12'b111101110000;
20'b01101101100100011111: color_data = 12'b111101110000;
20'b01101101100100100000: color_data = 12'b111101110000;
20'b01101101100100100100: color_data = 12'b111101110000;
20'b01101101100100100101: color_data = 12'b111101110000;
20'b01101101100100100110: color_data = 12'b111101110000;
20'b01101101100100100111: color_data = 12'b111101110000;
20'b01101101100100101000: color_data = 12'b111101110000;
20'b01101101100100101001: color_data = 12'b111101110000;
20'b01101101100100101010: color_data = 12'b111101110000;
20'b01101101100100101011: color_data = 12'b111101110000;
20'b01101101100100101100: color_data = 12'b111101110000;
20'b01101101100100101101: color_data = 12'b111101110000;
20'b01101101100100101110: color_data = 12'b111101110000;
20'b01101101100100101111: color_data = 12'b111101110000;
20'b01101101100100110000: color_data = 12'b111101110000;
20'b01101101100100110001: color_data = 12'b111101110000;
20'b01101101100100110010: color_data = 12'b111101110000;
20'b01101101100100110011: color_data = 12'b111101110000;
20'b01101101100100110100: color_data = 12'b111101110000;
20'b01101101100100110101: color_data = 12'b111101110000;
20'b01101101100100111001: color_data = 12'b111101110000;
20'b01101101100100111010: color_data = 12'b111101110000;
20'b01101101100100111011: color_data = 12'b111101110000;
20'b01101101100100111100: color_data = 12'b111101110000;
20'b01101101100100111101: color_data = 12'b111101110000;
20'b01101101100100111110: color_data = 12'b111101110000;
20'b01101101100100111111: color_data = 12'b111101110000;
20'b01101101100101000000: color_data = 12'b111101110000;
20'b01101101100101000001: color_data = 12'b111101110000;
20'b01101101100101000010: color_data = 12'b111101110000;
20'b01101101100101000011: color_data = 12'b111101110000;
20'b01101101100101000100: color_data = 12'b111101110000;
20'b01101101100101000101: color_data = 12'b111101110000;
20'b01101101100101000110: color_data = 12'b111101110000;
20'b01101101100101000111: color_data = 12'b111101110000;
20'b01101101100101001000: color_data = 12'b111101110000;
20'b01101101100101001001: color_data = 12'b111101110000;
20'b01101101100101001010: color_data = 12'b111101110000;
20'b01101101100101001110: color_data = 12'b000011110000;
20'b01101101100101001111: color_data = 12'b000011110000;
20'b01101101100101010000: color_data = 12'b000011110000;
20'b01101101100101010001: color_data = 12'b000011110000;
20'b01101101100101010010: color_data = 12'b000011110000;
20'b01101101100101010011: color_data = 12'b000011110000;
20'b01101101100101010100: color_data = 12'b000011110000;
20'b01101101100101010101: color_data = 12'b000011110000;
20'b01101101100101010110: color_data = 12'b000011110000;
20'b01101101100101010111: color_data = 12'b000011110000;
20'b01101101100101011000: color_data = 12'b000011110000;
20'b01101101100101011001: color_data = 12'b000011110000;
20'b01101101100101011010: color_data = 12'b000011110000;
20'b01101101100101011011: color_data = 12'b000011110000;
20'b01101101100101011100: color_data = 12'b000011110000;
20'b01101101100101011101: color_data = 12'b000011110000;
20'b01101101100101011110: color_data = 12'b000011110000;
20'b01101101100101011111: color_data = 12'b000011110000;
20'b01101101100101100011: color_data = 12'b111100001111;
20'b01101101100101100100: color_data = 12'b111100001111;
20'b01101101100101100101: color_data = 12'b111100001111;
20'b01101101100101100110: color_data = 12'b111100001111;
20'b01101101100101100111: color_data = 12'b111100001111;
20'b01101101100101101000: color_data = 12'b111100001111;
20'b01101101100101101001: color_data = 12'b111100001111;
20'b01101101100101101010: color_data = 12'b111100001111;
20'b01101101100101101011: color_data = 12'b111100001111;
20'b01101101100101101100: color_data = 12'b111100001111;
20'b01101101100101101101: color_data = 12'b111100001111;
20'b01101101100101101110: color_data = 12'b111100001111;
20'b01101101100101101111: color_data = 12'b111100001111;
20'b01101101100101110000: color_data = 12'b111100001111;
20'b01101101100101110001: color_data = 12'b111100001111;
20'b01101101100101110010: color_data = 12'b111100001111;
20'b01101101100101110011: color_data = 12'b111100001111;
20'b01101101100101110100: color_data = 12'b111100001111;
20'b01101101100101111000: color_data = 12'b111100000000;
20'b01101101100101111001: color_data = 12'b111100000000;
20'b01101101100101111010: color_data = 12'b111100000000;
20'b01101101100101111011: color_data = 12'b111100000000;
20'b01101101100101111100: color_data = 12'b111100000000;
20'b01101101100101111101: color_data = 12'b111100000000;
20'b01101101100101111110: color_data = 12'b111100000000;
20'b01101101100101111111: color_data = 12'b111100000000;
20'b01101101100110000000: color_data = 12'b111100000000;
20'b01101101100110000001: color_data = 12'b111100000000;
20'b01101101100110000010: color_data = 12'b111100000000;
20'b01101101100110000011: color_data = 12'b111100000000;
20'b01101101100110000100: color_data = 12'b111100000000;
20'b01101101100110000101: color_data = 12'b111100000000;
20'b01101101100110000110: color_data = 12'b111100000000;
20'b01101101100110000111: color_data = 12'b111100000000;
20'b01101101100110001000: color_data = 12'b111100000000;
20'b01101101100110001001: color_data = 12'b111100000000;
20'b01101101100110001101: color_data = 12'b111100000000;
20'b01101101100110001110: color_data = 12'b111100000000;
20'b01101101100110001111: color_data = 12'b111100000000;
20'b01101101100110010000: color_data = 12'b111100000000;
20'b01101101100110010001: color_data = 12'b111100000000;
20'b01101101100110010010: color_data = 12'b111100000000;
20'b01101101100110010011: color_data = 12'b111100000000;
20'b01101101100110010100: color_data = 12'b111100000000;
20'b01101101100110010101: color_data = 12'b111100000000;
20'b01101101100110010110: color_data = 12'b111100000000;
20'b01101101100110010111: color_data = 12'b111100000000;
20'b01101101100110011000: color_data = 12'b111100000000;
20'b01101101100110011001: color_data = 12'b111100000000;
20'b01101101100110011010: color_data = 12'b111100000000;
20'b01101101100110011011: color_data = 12'b111100000000;
20'b01101101100110011100: color_data = 12'b111100000000;
20'b01101101100110011101: color_data = 12'b111100000000;
20'b01101101100110011110: color_data = 12'b111100000000;
default: color_data = 12'b0;

	endcase
	end
endmodule