`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/29/2025 09:15:25 PM
// Design Name: 
// Module Name: game_over
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module game_over
	(
		input clk,
		input [9:0] row,
		input [9:0] col,
		output reg [11:0] color_data,
		input ce
	);
	    (* rom_style = "block" *)
	    
	reg [9:0] row_reg;
	reg [9:0] col_reg;
	always @(posedge clk)
		begin
		if (ce) begin
		row_reg <= row;
		col_reg <= col;
		end
		end
	always @(*) begin
	case ({row_reg, col_reg})
		20'b00010100100010100001: color_data = 12'b000011110111;
20'b00010100100010100010: color_data = 12'b000011110111;
20'b00010100100010100011: color_data = 12'b000011110111;
20'b00010100100010100100: color_data = 12'b000011110111;
20'b00010100100010100101: color_data = 12'b000011110111;
20'b00010100100010100110: color_data = 12'b000011110111;
20'b00010100100010100111: color_data = 12'b000011110111;
20'b00010100100010101000: color_data = 12'b000011110111;
20'b00010100100010101001: color_data = 12'b000011110111;
20'b00010100100010101010: color_data = 12'b000011110111;
20'b00010100100100001111: color_data = 12'b000000001111;
20'b00010100100100010000: color_data = 12'b000000001111;
20'b00010100100100010001: color_data = 12'b000000001111;
20'b00010100100100010010: color_data = 12'b000000001111;
20'b00010100100100010011: color_data = 12'b000000001111;
20'b00010100100100010100: color_data = 12'b000000001111;
20'b00010100100100010101: color_data = 12'b000000001111;
20'b00010100100100010110: color_data = 12'b000000001111;
20'b00010100100100010111: color_data = 12'b000000001111;
20'b00010100100100011000: color_data = 12'b000000001111;
20'b00010100100100011010: color_data = 12'b000000001111;
20'b00010100100100011011: color_data = 12'b000000001111;
20'b00010100100100011100: color_data = 12'b000000001111;
20'b00010100100100011101: color_data = 12'b000000001111;
20'b00010100100100011110: color_data = 12'b000000001111;
20'b00010100100100011111: color_data = 12'b000000001111;
20'b00010100100100100000: color_data = 12'b000000001111;
20'b00010100100100100001: color_data = 12'b000000001111;
20'b00010100100100100010: color_data = 12'b000000001111;
20'b00010100100100100011: color_data = 12'b000000001111;
20'b00010100110010100001: color_data = 12'b000011110111;
20'b00010100110010100010: color_data = 12'b000011110111;
20'b00010100110010100011: color_data = 12'b000011110111;
20'b00010100110010100100: color_data = 12'b000011110111;
20'b00010100110010100101: color_data = 12'b000011110111;
20'b00010100110010100110: color_data = 12'b000011110111;
20'b00010100110010100111: color_data = 12'b000011110111;
20'b00010100110010101000: color_data = 12'b000011110111;
20'b00010100110010101001: color_data = 12'b000011110111;
20'b00010100110010101010: color_data = 12'b000011110111;
20'b00010100110100001111: color_data = 12'b000000001111;
20'b00010100110100010000: color_data = 12'b000000001111;
20'b00010100110100010001: color_data = 12'b000000001111;
20'b00010100110100010010: color_data = 12'b000000001111;
20'b00010100110100010011: color_data = 12'b000000001111;
20'b00010100110100010100: color_data = 12'b000000001111;
20'b00010100110100010101: color_data = 12'b000000001111;
20'b00010100110100010110: color_data = 12'b000000001111;
20'b00010100110100010111: color_data = 12'b000000001111;
20'b00010100110100011000: color_data = 12'b000000001111;
20'b00010100110100011010: color_data = 12'b000000001111;
20'b00010100110100011011: color_data = 12'b000000001111;
20'b00010100110100011100: color_data = 12'b000000001111;
20'b00010100110100011101: color_data = 12'b000000001111;
20'b00010100110100011110: color_data = 12'b000000001111;
20'b00010100110100011111: color_data = 12'b000000001111;
20'b00010100110100100000: color_data = 12'b000000001111;
20'b00010100110100100001: color_data = 12'b000000001111;
20'b00010100110100100010: color_data = 12'b000000001111;
20'b00010100110100100011: color_data = 12'b000000001111;
20'b00010101000010100001: color_data = 12'b000011110111;
20'b00010101000010100010: color_data = 12'b000011110111;
20'b00010101000010100011: color_data = 12'b000011110111;
20'b00010101000010100100: color_data = 12'b000011110111;
20'b00010101000010100101: color_data = 12'b000011110111;
20'b00010101000010100110: color_data = 12'b000011110111;
20'b00010101000010100111: color_data = 12'b000011110111;
20'b00010101000010101000: color_data = 12'b000011110111;
20'b00010101000010101001: color_data = 12'b000011110111;
20'b00010101000010101010: color_data = 12'b000011110111;
20'b00010101000100001111: color_data = 12'b000000001111;
20'b00010101000100010000: color_data = 12'b000000001111;
20'b00010101000100010001: color_data = 12'b000000001111;
20'b00010101000100010010: color_data = 12'b000000001111;
20'b00010101000100010011: color_data = 12'b000000001111;
20'b00010101000100010100: color_data = 12'b000000001111;
20'b00010101000100010101: color_data = 12'b000000001111;
20'b00010101000100010110: color_data = 12'b000000001111;
20'b00010101000100010111: color_data = 12'b000000001111;
20'b00010101000100011000: color_data = 12'b000000001111;
20'b00010101000100011010: color_data = 12'b000000001111;
20'b00010101000100011011: color_data = 12'b000000001111;
20'b00010101000100011100: color_data = 12'b000000001111;
20'b00010101000100011101: color_data = 12'b000000001111;
20'b00010101000100011110: color_data = 12'b000000001111;
20'b00010101000100011111: color_data = 12'b000000001111;
20'b00010101000100100000: color_data = 12'b000000001111;
20'b00010101000100100001: color_data = 12'b000000001111;
20'b00010101000100100010: color_data = 12'b000000001111;
20'b00010101000100100011: color_data = 12'b000000001111;
20'b00010101010010100001: color_data = 12'b000011110111;
20'b00010101010010100010: color_data = 12'b000011110111;
20'b00010101010010100011: color_data = 12'b000011110111;
20'b00010101010010100100: color_data = 12'b000011110111;
20'b00010101010010100101: color_data = 12'b000011110111;
20'b00010101010010100110: color_data = 12'b000011110111;
20'b00010101010010100111: color_data = 12'b000011110111;
20'b00010101010010101000: color_data = 12'b000011110111;
20'b00010101010010101001: color_data = 12'b000011110111;
20'b00010101010010101010: color_data = 12'b000011110111;
20'b00010101010100001111: color_data = 12'b000000001111;
20'b00010101010100010000: color_data = 12'b000000001111;
20'b00010101010100010001: color_data = 12'b000000001111;
20'b00010101010100010010: color_data = 12'b000000001111;
20'b00010101010100010011: color_data = 12'b000000001111;
20'b00010101010100010100: color_data = 12'b000000001111;
20'b00010101010100010101: color_data = 12'b000000001111;
20'b00010101010100010110: color_data = 12'b000000001111;
20'b00010101010100010111: color_data = 12'b000000001111;
20'b00010101010100011000: color_data = 12'b000000001111;
20'b00010101010100011010: color_data = 12'b000000001111;
20'b00010101010100011011: color_data = 12'b000000001111;
20'b00010101010100011100: color_data = 12'b000000001111;
20'b00010101010100011101: color_data = 12'b000000001111;
20'b00010101010100011110: color_data = 12'b000000001111;
20'b00010101010100011111: color_data = 12'b000000001111;
20'b00010101010100100000: color_data = 12'b000000001111;
20'b00010101010100100001: color_data = 12'b000000001111;
20'b00010101010100100010: color_data = 12'b000000001111;
20'b00010101010100100011: color_data = 12'b000000001111;
20'b00010101100010100001: color_data = 12'b000011110111;
20'b00010101100010100010: color_data = 12'b000011110111;
20'b00010101100010100011: color_data = 12'b000011110111;
20'b00010101100010100100: color_data = 12'b000011110111;
20'b00010101100010100101: color_data = 12'b000011110111;
20'b00010101100010100110: color_data = 12'b000011110111;
20'b00010101100010100111: color_data = 12'b000011110111;
20'b00010101100010101000: color_data = 12'b000011110111;
20'b00010101100010101001: color_data = 12'b000011110111;
20'b00010101100010101010: color_data = 12'b000011110111;
20'b00010101100100001111: color_data = 12'b000000001111;
20'b00010101100100010000: color_data = 12'b000000001111;
20'b00010101100100010001: color_data = 12'b000000001111;
20'b00010101100100010010: color_data = 12'b000000001111;
20'b00010101100100010011: color_data = 12'b000000001111;
20'b00010101100100010100: color_data = 12'b000000001111;
20'b00010101100100010101: color_data = 12'b000000001111;
20'b00010101100100010110: color_data = 12'b000000001111;
20'b00010101100100010111: color_data = 12'b000000001111;
20'b00010101100100011000: color_data = 12'b000000001111;
20'b00010101100100011010: color_data = 12'b000000001111;
20'b00010101100100011011: color_data = 12'b000000001111;
20'b00010101100100011100: color_data = 12'b000000001111;
20'b00010101100100011101: color_data = 12'b000000001111;
20'b00010101100100011110: color_data = 12'b000000001111;
20'b00010101100100011111: color_data = 12'b000000001111;
20'b00010101100100100000: color_data = 12'b000000001111;
20'b00010101100100100001: color_data = 12'b000000001111;
20'b00010101100100100010: color_data = 12'b000000001111;
20'b00010101100100100011: color_data = 12'b000000001111;
20'b00010101110010100001: color_data = 12'b000011110111;
20'b00010101110010100010: color_data = 12'b000011110111;
20'b00010101110010100011: color_data = 12'b000011110111;
20'b00010101110010100100: color_data = 12'b000011110111;
20'b00010101110010100101: color_data = 12'b000011110111;
20'b00010101110010100110: color_data = 12'b000011110111;
20'b00010101110010100111: color_data = 12'b000011110111;
20'b00010101110010101000: color_data = 12'b000011110111;
20'b00010101110010101001: color_data = 12'b000011110111;
20'b00010101110010101010: color_data = 12'b000011110111;
20'b00010101110100001111: color_data = 12'b000000001111;
20'b00010101110100010000: color_data = 12'b000000001111;
20'b00010101110100010001: color_data = 12'b000000001111;
20'b00010101110100010010: color_data = 12'b000000001111;
20'b00010101110100010011: color_data = 12'b000000001111;
20'b00010101110100010100: color_data = 12'b000000001111;
20'b00010101110100010101: color_data = 12'b000000001111;
20'b00010101110100010110: color_data = 12'b000000001111;
20'b00010101110100010111: color_data = 12'b000000001111;
20'b00010101110100011000: color_data = 12'b000000001111;
20'b00010101110100011010: color_data = 12'b000000001111;
20'b00010101110100011011: color_data = 12'b000000001111;
20'b00010101110100011100: color_data = 12'b000000001111;
20'b00010101110100011101: color_data = 12'b000000001111;
20'b00010101110100011110: color_data = 12'b000000001111;
20'b00010101110100011111: color_data = 12'b000000001111;
20'b00010101110100100000: color_data = 12'b000000001111;
20'b00010101110100100001: color_data = 12'b000000001111;
20'b00010101110100100010: color_data = 12'b000000001111;
20'b00010101110100100011: color_data = 12'b000000001111;
20'b00010101110110011110: color_data = 12'b000011110111;
20'b00010101110110011111: color_data = 12'b000011110111;
20'b00010101110110100000: color_data = 12'b000011110111;
20'b00010101110110100001: color_data = 12'b000011110111;
20'b00010101110110100010: color_data = 12'b000011110111;
20'b00010101110110100011: color_data = 12'b000011110111;
20'b00010101110110100100: color_data = 12'b000011110111;
20'b00010101110110100101: color_data = 12'b000011110111;
20'b00010101110110100110: color_data = 12'b000011110111;
20'b00010101110110100111: color_data = 12'b000011110111;
20'b00010101110110101001: color_data = 12'b000011110111;
20'b00010101110110101010: color_data = 12'b000011110111;
20'b00010101110110101011: color_data = 12'b000011110111;
20'b00010101110110101100: color_data = 12'b000011110111;
20'b00010101110110101101: color_data = 12'b000011110111;
20'b00010101110110101110: color_data = 12'b000011110111;
20'b00010101110110101111: color_data = 12'b000011110111;
20'b00010101110110110000: color_data = 12'b000011110111;
20'b00010101110110110001: color_data = 12'b000011110111;
20'b00010101110110110010: color_data = 12'b000011110111;
20'b00010110000010100001: color_data = 12'b000011110111;
20'b00010110000010100010: color_data = 12'b000011110111;
20'b00010110000010100011: color_data = 12'b000011110111;
20'b00010110000010100100: color_data = 12'b000011110111;
20'b00010110000010100101: color_data = 12'b000011110111;
20'b00010110000010100110: color_data = 12'b000011110111;
20'b00010110000010100111: color_data = 12'b000011110111;
20'b00010110000010101000: color_data = 12'b000011110111;
20'b00010110000010101001: color_data = 12'b000011110111;
20'b00010110000010101010: color_data = 12'b000011110111;
20'b00010110000100001111: color_data = 12'b000000001111;
20'b00010110000100010000: color_data = 12'b000000001111;
20'b00010110000100010001: color_data = 12'b000000001111;
20'b00010110000100010010: color_data = 12'b000000001111;
20'b00010110000100010011: color_data = 12'b000000001111;
20'b00010110000100010100: color_data = 12'b000000001111;
20'b00010110000100010101: color_data = 12'b000000001111;
20'b00010110000100010110: color_data = 12'b000000001111;
20'b00010110000100010111: color_data = 12'b000000001111;
20'b00010110000100011000: color_data = 12'b000000001111;
20'b00010110000100011010: color_data = 12'b000000001111;
20'b00010110000100011011: color_data = 12'b000000001111;
20'b00010110000100011100: color_data = 12'b000000001111;
20'b00010110000100011101: color_data = 12'b000000001111;
20'b00010110000100011110: color_data = 12'b000000001111;
20'b00010110000100011111: color_data = 12'b000000001111;
20'b00010110000100100000: color_data = 12'b000000001111;
20'b00010110000100100001: color_data = 12'b000000001111;
20'b00010110000100100010: color_data = 12'b000000001111;
20'b00010110000100100011: color_data = 12'b000000001111;
20'b00010110000110011110: color_data = 12'b000011110111;
20'b00010110000110011111: color_data = 12'b000011110111;
20'b00010110000110100000: color_data = 12'b000011110111;
20'b00010110000110100001: color_data = 12'b000011110111;
20'b00010110000110100010: color_data = 12'b000011110111;
20'b00010110000110100011: color_data = 12'b000011110111;
20'b00010110000110100100: color_data = 12'b000011110111;
20'b00010110000110100101: color_data = 12'b000011110111;
20'b00010110000110100110: color_data = 12'b000011110111;
20'b00010110000110100111: color_data = 12'b000011110111;
20'b00010110000110101001: color_data = 12'b000011110111;
20'b00010110000110101010: color_data = 12'b000011110111;
20'b00010110000110101011: color_data = 12'b000011110111;
20'b00010110000110101100: color_data = 12'b000011110111;
20'b00010110000110101101: color_data = 12'b000011110111;
20'b00010110000110101110: color_data = 12'b000011110111;
20'b00010110000110101111: color_data = 12'b000011110111;
20'b00010110000110110000: color_data = 12'b000011110111;
20'b00010110000110110001: color_data = 12'b000011110111;
20'b00010110000110110010: color_data = 12'b000011110111;
20'b00010110010010100001: color_data = 12'b000011110111;
20'b00010110010010100010: color_data = 12'b000011110111;
20'b00010110010010100011: color_data = 12'b000011110111;
20'b00010110010010100100: color_data = 12'b000011110111;
20'b00010110010010100101: color_data = 12'b000011110111;
20'b00010110010010100110: color_data = 12'b000011110111;
20'b00010110010010100111: color_data = 12'b000011110111;
20'b00010110010010101000: color_data = 12'b000011110111;
20'b00010110010010101001: color_data = 12'b000011110111;
20'b00010110010010101010: color_data = 12'b000011110111;
20'b00010110010100001111: color_data = 12'b000000001111;
20'b00010110010100010000: color_data = 12'b000000001111;
20'b00010110010100010001: color_data = 12'b000000001111;
20'b00010110010100010010: color_data = 12'b000000001111;
20'b00010110010100010011: color_data = 12'b000000001111;
20'b00010110010100010100: color_data = 12'b000000001111;
20'b00010110010100010101: color_data = 12'b000000001111;
20'b00010110010100010110: color_data = 12'b000000001111;
20'b00010110010100010111: color_data = 12'b000000001111;
20'b00010110010100011000: color_data = 12'b000000001111;
20'b00010110010100011010: color_data = 12'b000000001111;
20'b00010110010100011011: color_data = 12'b000000001111;
20'b00010110010100011100: color_data = 12'b000000001111;
20'b00010110010100011101: color_data = 12'b000000001111;
20'b00010110010100011110: color_data = 12'b000000001111;
20'b00010110010100011111: color_data = 12'b000000001111;
20'b00010110010100100000: color_data = 12'b000000001111;
20'b00010110010100100001: color_data = 12'b000000001111;
20'b00010110010100100010: color_data = 12'b000000001111;
20'b00010110010100100011: color_data = 12'b000000001111;
20'b00010110010110011110: color_data = 12'b000011110111;
20'b00010110010110011111: color_data = 12'b000011110111;
20'b00010110010110100000: color_data = 12'b000011110111;
20'b00010110010110100001: color_data = 12'b000011110111;
20'b00010110010110100010: color_data = 12'b000011110111;
20'b00010110010110100011: color_data = 12'b000011110111;
20'b00010110010110100100: color_data = 12'b000011110111;
20'b00010110010110100101: color_data = 12'b000011110111;
20'b00010110010110100110: color_data = 12'b000011110111;
20'b00010110010110100111: color_data = 12'b000011110111;
20'b00010110010110101001: color_data = 12'b000011110111;
20'b00010110010110101010: color_data = 12'b000011110111;
20'b00010110010110101011: color_data = 12'b000011110111;
20'b00010110010110101100: color_data = 12'b000011110111;
20'b00010110010110101101: color_data = 12'b000011110111;
20'b00010110010110101110: color_data = 12'b000011110111;
20'b00010110010110101111: color_data = 12'b000011110111;
20'b00010110010110110000: color_data = 12'b000011110111;
20'b00010110010110110001: color_data = 12'b000011110111;
20'b00010110010110110010: color_data = 12'b000011110111;
20'b00010110100010100001: color_data = 12'b000011110111;
20'b00010110100010100010: color_data = 12'b000011110111;
20'b00010110100010100011: color_data = 12'b000011110111;
20'b00010110100010100100: color_data = 12'b000011110111;
20'b00010110100010100101: color_data = 12'b000011110111;
20'b00010110100010100110: color_data = 12'b000011110111;
20'b00010110100010100111: color_data = 12'b000011110111;
20'b00010110100010101000: color_data = 12'b000011110111;
20'b00010110100010101001: color_data = 12'b000011110111;
20'b00010110100010101010: color_data = 12'b000011110111;
20'b00010110100100001111: color_data = 12'b000000001111;
20'b00010110100100010000: color_data = 12'b000000001111;
20'b00010110100100010001: color_data = 12'b000000001111;
20'b00010110100100010010: color_data = 12'b000000001111;
20'b00010110100100010011: color_data = 12'b000000001111;
20'b00010110100100010100: color_data = 12'b000000001111;
20'b00010110100100010101: color_data = 12'b000000001111;
20'b00010110100100010110: color_data = 12'b000000001111;
20'b00010110100100010111: color_data = 12'b000000001111;
20'b00010110100100011000: color_data = 12'b000000001111;
20'b00010110100100011010: color_data = 12'b000000001111;
20'b00010110100100011011: color_data = 12'b000000001111;
20'b00010110100100011100: color_data = 12'b000000001111;
20'b00010110100100011101: color_data = 12'b000000001111;
20'b00010110100100011110: color_data = 12'b000000001111;
20'b00010110100100011111: color_data = 12'b000000001111;
20'b00010110100100100000: color_data = 12'b000000001111;
20'b00010110100100100001: color_data = 12'b000000001111;
20'b00010110100100100010: color_data = 12'b000000001111;
20'b00010110100100100011: color_data = 12'b000000001111;
20'b00010110100110011110: color_data = 12'b000011110111;
20'b00010110100110011111: color_data = 12'b000011110111;
20'b00010110100110100000: color_data = 12'b000011110111;
20'b00010110100110100001: color_data = 12'b000011110111;
20'b00010110100110100010: color_data = 12'b000011110111;
20'b00010110100110100011: color_data = 12'b000011110111;
20'b00010110100110100100: color_data = 12'b000011110111;
20'b00010110100110100101: color_data = 12'b000011110111;
20'b00010110100110100110: color_data = 12'b000011110111;
20'b00010110100110100111: color_data = 12'b000011110111;
20'b00010110100110101001: color_data = 12'b000011110111;
20'b00010110100110101010: color_data = 12'b000011110111;
20'b00010110100110101011: color_data = 12'b000011110111;
20'b00010110100110101100: color_data = 12'b000011110111;
20'b00010110100110101101: color_data = 12'b000011110111;
20'b00010110100110101110: color_data = 12'b000011110111;
20'b00010110100110101111: color_data = 12'b000011110111;
20'b00010110100110110000: color_data = 12'b000011110111;
20'b00010110100110110001: color_data = 12'b000011110111;
20'b00010110100110110010: color_data = 12'b000011110111;
20'b00010110110010100001: color_data = 12'b000011110111;
20'b00010110110010100010: color_data = 12'b000011110111;
20'b00010110110010100011: color_data = 12'b000011110111;
20'b00010110110010100100: color_data = 12'b000011110111;
20'b00010110110010100101: color_data = 12'b000011110111;
20'b00010110110010100110: color_data = 12'b000011110111;
20'b00010110110010100111: color_data = 12'b000011110111;
20'b00010110110010101000: color_data = 12'b000011110111;
20'b00010110110010101001: color_data = 12'b000011110111;
20'b00010110110010101010: color_data = 12'b000011110111;
20'b00010110110100001111: color_data = 12'b000000001111;
20'b00010110110100010000: color_data = 12'b000000001111;
20'b00010110110100010001: color_data = 12'b000000001111;
20'b00010110110100010010: color_data = 12'b000000001111;
20'b00010110110100010011: color_data = 12'b000000001111;
20'b00010110110100010100: color_data = 12'b000000001111;
20'b00010110110100010101: color_data = 12'b000000001111;
20'b00010110110100010110: color_data = 12'b000000001111;
20'b00010110110100010111: color_data = 12'b000000001111;
20'b00010110110100011000: color_data = 12'b000000001111;
20'b00010110110100011010: color_data = 12'b000000001111;
20'b00010110110100011011: color_data = 12'b000000001111;
20'b00010110110100011100: color_data = 12'b000000001111;
20'b00010110110100011101: color_data = 12'b000000001111;
20'b00010110110100011110: color_data = 12'b000000001111;
20'b00010110110100011111: color_data = 12'b000000001111;
20'b00010110110100100000: color_data = 12'b000000001111;
20'b00010110110100100001: color_data = 12'b000000001111;
20'b00010110110100100010: color_data = 12'b000000001111;
20'b00010110110100100011: color_data = 12'b000000001111;
20'b00010110110110011110: color_data = 12'b000011110111;
20'b00010110110110011111: color_data = 12'b000011110111;
20'b00010110110110100000: color_data = 12'b000011110111;
20'b00010110110110100001: color_data = 12'b000011110111;
20'b00010110110110100010: color_data = 12'b000011110111;
20'b00010110110110100011: color_data = 12'b000011110111;
20'b00010110110110100100: color_data = 12'b000011110111;
20'b00010110110110100101: color_data = 12'b000011110111;
20'b00010110110110100110: color_data = 12'b000011110111;
20'b00010110110110100111: color_data = 12'b000011110111;
20'b00010110110110101001: color_data = 12'b000011110111;
20'b00010110110110101010: color_data = 12'b000011110111;
20'b00010110110110101011: color_data = 12'b000011110111;
20'b00010110110110101100: color_data = 12'b000011110111;
20'b00010110110110101101: color_data = 12'b000011110111;
20'b00010110110110101110: color_data = 12'b000011110111;
20'b00010110110110101111: color_data = 12'b000011110111;
20'b00010110110110110000: color_data = 12'b000011110111;
20'b00010110110110110001: color_data = 12'b000011110111;
20'b00010110110110110010: color_data = 12'b000011110111;
20'b00010111000110011110: color_data = 12'b000011110111;
20'b00010111000110011111: color_data = 12'b000011110111;
20'b00010111000110100000: color_data = 12'b000011110111;
20'b00010111000110100001: color_data = 12'b000011110111;
20'b00010111000110100010: color_data = 12'b000011110111;
20'b00010111000110100011: color_data = 12'b000011110111;
20'b00010111000110100100: color_data = 12'b000011110111;
20'b00010111000110100101: color_data = 12'b000011110111;
20'b00010111000110100110: color_data = 12'b000011110111;
20'b00010111000110100111: color_data = 12'b000011110111;
20'b00010111000110101001: color_data = 12'b000011110111;
20'b00010111000110101010: color_data = 12'b000011110111;
20'b00010111000110101011: color_data = 12'b000011110111;
20'b00010111000110101100: color_data = 12'b000011110111;
20'b00010111000110101101: color_data = 12'b000011110111;
20'b00010111000110101110: color_data = 12'b000011110111;
20'b00010111000110101111: color_data = 12'b000011110111;
20'b00010111000110110000: color_data = 12'b000011110111;
20'b00010111000110110001: color_data = 12'b000011110111;
20'b00010111000110110010: color_data = 12'b000011110111;
20'b00010111010010010110: color_data = 12'b000011110111;
20'b00010111010010010111: color_data = 12'b000011110111;
20'b00010111010010011000: color_data = 12'b000011110111;
20'b00010111010010011001: color_data = 12'b000011110111;
20'b00010111010010011010: color_data = 12'b000011110111;
20'b00010111010010011011: color_data = 12'b000011110111;
20'b00010111010010011100: color_data = 12'b000011110111;
20'b00010111010010011101: color_data = 12'b000011110111;
20'b00010111010010011110: color_data = 12'b000011110111;
20'b00010111010010011111: color_data = 12'b000011110111;
20'b00010111010010100001: color_data = 12'b000011110111;
20'b00010111010010100010: color_data = 12'b000011110111;
20'b00010111010010100011: color_data = 12'b000011110111;
20'b00010111010010100100: color_data = 12'b000011110111;
20'b00010111010010100101: color_data = 12'b000011110111;
20'b00010111010010100110: color_data = 12'b000011110111;
20'b00010111010010100111: color_data = 12'b000011110111;
20'b00010111010010101000: color_data = 12'b000011110111;
20'b00010111010010101001: color_data = 12'b000011110111;
20'b00010111010010101010: color_data = 12'b000011110111;
20'b00010111010100011010: color_data = 12'b000000001111;
20'b00010111010100011011: color_data = 12'b000000001111;
20'b00010111010100011100: color_data = 12'b000000001111;
20'b00010111010100011101: color_data = 12'b000000001111;
20'b00010111010100011110: color_data = 12'b000000001111;
20'b00010111010100011111: color_data = 12'b000000001111;
20'b00010111010100100000: color_data = 12'b000000001111;
20'b00010111010100100001: color_data = 12'b000000001111;
20'b00010111010100100010: color_data = 12'b000000001111;
20'b00010111010100100011: color_data = 12'b000000001111;
20'b00010111010110011110: color_data = 12'b000011110111;
20'b00010111010110011111: color_data = 12'b000011110111;
20'b00010111010110100000: color_data = 12'b000011110111;
20'b00010111010110100001: color_data = 12'b000011110111;
20'b00010111010110100010: color_data = 12'b000011110111;
20'b00010111010110100011: color_data = 12'b000011110111;
20'b00010111010110100100: color_data = 12'b000011110111;
20'b00010111010110100101: color_data = 12'b000011110111;
20'b00010111010110100110: color_data = 12'b000011110111;
20'b00010111010110100111: color_data = 12'b000011110111;
20'b00010111010110101001: color_data = 12'b000011110111;
20'b00010111010110101010: color_data = 12'b000011110111;
20'b00010111010110101011: color_data = 12'b000011110111;
20'b00010111010110101100: color_data = 12'b000011110111;
20'b00010111010110101101: color_data = 12'b000011110111;
20'b00010111010110101110: color_data = 12'b000011110111;
20'b00010111010110101111: color_data = 12'b000011110111;
20'b00010111010110110000: color_data = 12'b000011110111;
20'b00010111010110110001: color_data = 12'b000011110111;
20'b00010111010110110010: color_data = 12'b000011110111;
20'b00010111100010010110: color_data = 12'b000011110111;
20'b00010111100010010111: color_data = 12'b000011110111;
20'b00010111100010011000: color_data = 12'b000011110111;
20'b00010111100010011001: color_data = 12'b000011110111;
20'b00010111100010011010: color_data = 12'b000011110111;
20'b00010111100010011011: color_data = 12'b000011110111;
20'b00010111100010011100: color_data = 12'b000011110111;
20'b00010111100010011101: color_data = 12'b000011110111;
20'b00010111100010011110: color_data = 12'b000011110111;
20'b00010111100010011111: color_data = 12'b000011110111;
20'b00010111100010100001: color_data = 12'b000011110111;
20'b00010111100010100010: color_data = 12'b000011110111;
20'b00010111100010100011: color_data = 12'b000011110111;
20'b00010111100010100100: color_data = 12'b000011110111;
20'b00010111100010100101: color_data = 12'b000011110111;
20'b00010111100010100110: color_data = 12'b000011110111;
20'b00010111100010100111: color_data = 12'b000011110111;
20'b00010111100010101000: color_data = 12'b000011110111;
20'b00010111100010101001: color_data = 12'b000011110111;
20'b00010111100010101010: color_data = 12'b000011110111;
20'b00010111100100011010: color_data = 12'b000000001111;
20'b00010111100100011011: color_data = 12'b000000001111;
20'b00010111100100011100: color_data = 12'b000000001111;
20'b00010111100100011101: color_data = 12'b000000001111;
20'b00010111100100011110: color_data = 12'b000000001111;
20'b00010111100100011111: color_data = 12'b000000001111;
20'b00010111100100100000: color_data = 12'b000000001111;
20'b00010111100100100001: color_data = 12'b000000001111;
20'b00010111100100100010: color_data = 12'b000000001111;
20'b00010111100100100011: color_data = 12'b000000001111;
20'b00010111100110011110: color_data = 12'b000011110111;
20'b00010111100110011111: color_data = 12'b000011110111;
20'b00010111100110100000: color_data = 12'b000011110111;
20'b00010111100110100001: color_data = 12'b000011110111;
20'b00010111100110100010: color_data = 12'b000011110111;
20'b00010111100110100011: color_data = 12'b000011110111;
20'b00010111100110100100: color_data = 12'b000011110111;
20'b00010111100110100101: color_data = 12'b000011110111;
20'b00010111100110100110: color_data = 12'b000011110111;
20'b00010111100110100111: color_data = 12'b000011110111;
20'b00010111100110101001: color_data = 12'b000011110111;
20'b00010111100110101010: color_data = 12'b000011110111;
20'b00010111100110101011: color_data = 12'b000011110111;
20'b00010111100110101100: color_data = 12'b000011110111;
20'b00010111100110101101: color_data = 12'b000011110111;
20'b00010111100110101110: color_data = 12'b000011110111;
20'b00010111100110101111: color_data = 12'b000011110111;
20'b00010111100110110000: color_data = 12'b000011110111;
20'b00010111100110110001: color_data = 12'b000011110111;
20'b00010111100110110010: color_data = 12'b000011110111;
20'b00010111110010010110: color_data = 12'b000011110111;
20'b00010111110010010111: color_data = 12'b000011110111;
20'b00010111110010011000: color_data = 12'b000011110111;
20'b00010111110010011001: color_data = 12'b000011110111;
20'b00010111110010011010: color_data = 12'b000011110111;
20'b00010111110010011011: color_data = 12'b000011110111;
20'b00010111110010011100: color_data = 12'b000011110111;
20'b00010111110010011101: color_data = 12'b000011110111;
20'b00010111110010011110: color_data = 12'b000011110111;
20'b00010111110010011111: color_data = 12'b000011110111;
20'b00010111110010100001: color_data = 12'b000011110111;
20'b00010111110010100010: color_data = 12'b000011110111;
20'b00010111110010100011: color_data = 12'b000011110111;
20'b00010111110010100100: color_data = 12'b000011110111;
20'b00010111110010100101: color_data = 12'b000011110111;
20'b00010111110010100110: color_data = 12'b000011110111;
20'b00010111110010100111: color_data = 12'b000011110111;
20'b00010111110010101000: color_data = 12'b000011110111;
20'b00010111110010101001: color_data = 12'b000011110111;
20'b00010111110010101010: color_data = 12'b000011110111;
20'b00010111110100011010: color_data = 12'b000000001111;
20'b00010111110100011011: color_data = 12'b000000001111;
20'b00010111110100011100: color_data = 12'b000000001111;
20'b00010111110100011101: color_data = 12'b000000001111;
20'b00010111110100011110: color_data = 12'b000000001111;
20'b00010111110100011111: color_data = 12'b000000001111;
20'b00010111110100100000: color_data = 12'b000000001111;
20'b00010111110100100001: color_data = 12'b000000001111;
20'b00010111110100100010: color_data = 12'b000000001111;
20'b00010111110100100011: color_data = 12'b000000001111;
20'b00010111110110011110: color_data = 12'b000011110111;
20'b00010111110110011111: color_data = 12'b000011110111;
20'b00010111110110100000: color_data = 12'b000011110111;
20'b00010111110110100001: color_data = 12'b000011110111;
20'b00010111110110100010: color_data = 12'b000011110111;
20'b00010111110110100011: color_data = 12'b000011110111;
20'b00010111110110100100: color_data = 12'b000011110111;
20'b00010111110110100101: color_data = 12'b000011110111;
20'b00010111110110100110: color_data = 12'b000011110111;
20'b00010111110110100111: color_data = 12'b000011110111;
20'b00010111110110101001: color_data = 12'b000011110111;
20'b00010111110110101010: color_data = 12'b000011110111;
20'b00010111110110101011: color_data = 12'b000011110111;
20'b00010111110110101100: color_data = 12'b000011110111;
20'b00010111110110101101: color_data = 12'b000011110111;
20'b00010111110110101110: color_data = 12'b000011110111;
20'b00010111110110101111: color_data = 12'b000011110111;
20'b00010111110110110000: color_data = 12'b000011110111;
20'b00010111110110110001: color_data = 12'b000011110111;
20'b00010111110110110010: color_data = 12'b000011110111;
20'b00011000000010010110: color_data = 12'b000011110111;
20'b00011000000010010111: color_data = 12'b000011110111;
20'b00011000000010011000: color_data = 12'b000011110111;
20'b00011000000010011001: color_data = 12'b000011110111;
20'b00011000000010011010: color_data = 12'b000011110111;
20'b00011000000010011011: color_data = 12'b000011110111;
20'b00011000000010011100: color_data = 12'b000011110111;
20'b00011000000010011101: color_data = 12'b000011110111;
20'b00011000000010011110: color_data = 12'b000011110111;
20'b00011000000010011111: color_data = 12'b000011110111;
20'b00011000000010100001: color_data = 12'b000011110111;
20'b00011000000010100010: color_data = 12'b000011110111;
20'b00011000000010100011: color_data = 12'b000011110111;
20'b00011000000010100100: color_data = 12'b000011110111;
20'b00011000000010100101: color_data = 12'b000011110111;
20'b00011000000010100110: color_data = 12'b000011110111;
20'b00011000000010100111: color_data = 12'b000011110111;
20'b00011000000010101000: color_data = 12'b000011110111;
20'b00011000000010101001: color_data = 12'b000011110111;
20'b00011000000010101010: color_data = 12'b000011110111;
20'b00011000000100011010: color_data = 12'b000000001111;
20'b00011000000100011011: color_data = 12'b000000001111;
20'b00011000000100011100: color_data = 12'b000000001111;
20'b00011000000100011101: color_data = 12'b000000001111;
20'b00011000000100011110: color_data = 12'b000000001111;
20'b00011000000100011111: color_data = 12'b000000001111;
20'b00011000000100100000: color_data = 12'b000000001111;
20'b00011000000100100001: color_data = 12'b000000001111;
20'b00011000000100100010: color_data = 12'b000000001111;
20'b00011000000100100011: color_data = 12'b000000001111;
20'b00011000010010010110: color_data = 12'b000011110111;
20'b00011000010010010111: color_data = 12'b000011110111;
20'b00011000010010011000: color_data = 12'b000011110111;
20'b00011000010010011001: color_data = 12'b000011110111;
20'b00011000010010011010: color_data = 12'b000011110111;
20'b00011000010010011011: color_data = 12'b000011110111;
20'b00011000010010011100: color_data = 12'b000011110111;
20'b00011000010010011101: color_data = 12'b000011110111;
20'b00011000010010011110: color_data = 12'b000011110111;
20'b00011000010010011111: color_data = 12'b000011110111;
20'b00011000010010100001: color_data = 12'b000011110111;
20'b00011000010010100010: color_data = 12'b000011110111;
20'b00011000010010100011: color_data = 12'b000011110111;
20'b00011000010010100100: color_data = 12'b000011110111;
20'b00011000010010100101: color_data = 12'b000011110111;
20'b00011000010010100110: color_data = 12'b000011110111;
20'b00011000010010100111: color_data = 12'b000011110111;
20'b00011000010010101000: color_data = 12'b000011110111;
20'b00011000010010101001: color_data = 12'b000011110111;
20'b00011000010010101010: color_data = 12'b000011110111;
20'b00011000010100011010: color_data = 12'b000000001111;
20'b00011000010100011011: color_data = 12'b000000001111;
20'b00011000010100011100: color_data = 12'b000000001111;
20'b00011000010100011101: color_data = 12'b000000001111;
20'b00011000010100011110: color_data = 12'b000000001111;
20'b00011000010100011111: color_data = 12'b000000001111;
20'b00011000010100100000: color_data = 12'b000000001111;
20'b00011000010100100001: color_data = 12'b000000001111;
20'b00011000010100100010: color_data = 12'b000000001111;
20'b00011000010100100011: color_data = 12'b000000001111;
20'b00011000010110011110: color_data = 12'b000011110111;
20'b00011000010110011111: color_data = 12'b000011110111;
20'b00011000010110100000: color_data = 12'b000011110111;
20'b00011000010110100001: color_data = 12'b000011110111;
20'b00011000010110100010: color_data = 12'b000011110111;
20'b00011000010110100011: color_data = 12'b000011110111;
20'b00011000010110100100: color_data = 12'b000011110111;
20'b00011000010110100101: color_data = 12'b000011110111;
20'b00011000010110100110: color_data = 12'b000011110111;
20'b00011000010110100111: color_data = 12'b000011110111;
20'b00011000100010010110: color_data = 12'b000011110111;
20'b00011000100010010111: color_data = 12'b000011110111;
20'b00011000100010011000: color_data = 12'b000011110111;
20'b00011000100010011001: color_data = 12'b000011110111;
20'b00011000100010011010: color_data = 12'b000011110111;
20'b00011000100010011011: color_data = 12'b000011110111;
20'b00011000100010011100: color_data = 12'b000011110111;
20'b00011000100010011101: color_data = 12'b000011110111;
20'b00011000100010011110: color_data = 12'b000011110111;
20'b00011000100010011111: color_data = 12'b000011110111;
20'b00011000100010100001: color_data = 12'b000011110111;
20'b00011000100010100010: color_data = 12'b000011110111;
20'b00011000100010100011: color_data = 12'b000011110111;
20'b00011000100010100100: color_data = 12'b000011110111;
20'b00011000100010100101: color_data = 12'b000011110111;
20'b00011000100010100110: color_data = 12'b000011110111;
20'b00011000100010100111: color_data = 12'b000011110111;
20'b00011000100010101000: color_data = 12'b000011110111;
20'b00011000100010101001: color_data = 12'b000011110111;
20'b00011000100010101010: color_data = 12'b000011110111;
20'b00011000100100011010: color_data = 12'b000000001111;
20'b00011000100100011011: color_data = 12'b000000001111;
20'b00011000100100011100: color_data = 12'b000000001111;
20'b00011000100100011101: color_data = 12'b000000001111;
20'b00011000100100011110: color_data = 12'b000000001111;
20'b00011000100100011111: color_data = 12'b000000001111;
20'b00011000100100100000: color_data = 12'b000000001111;
20'b00011000100100100001: color_data = 12'b000000001111;
20'b00011000100100100010: color_data = 12'b000000001111;
20'b00011000100100100011: color_data = 12'b000000001111;
20'b00011000100110011110: color_data = 12'b000011110111;
20'b00011000100110011111: color_data = 12'b000011110111;
20'b00011000100110100000: color_data = 12'b000011110111;
20'b00011000100110100001: color_data = 12'b000011110111;
20'b00011000100110100010: color_data = 12'b000011110111;
20'b00011000100110100011: color_data = 12'b000011110111;
20'b00011000100110100100: color_data = 12'b000011110111;
20'b00011000100110100101: color_data = 12'b000011110111;
20'b00011000100110100110: color_data = 12'b000011110111;
20'b00011000100110100111: color_data = 12'b000011110111;
20'b00011000110010010110: color_data = 12'b000011110111;
20'b00011000110010010111: color_data = 12'b000011110111;
20'b00011000110010011000: color_data = 12'b000011110111;
20'b00011000110010011001: color_data = 12'b000011110111;
20'b00011000110010011010: color_data = 12'b000011110111;
20'b00011000110010011011: color_data = 12'b000011110111;
20'b00011000110010011100: color_data = 12'b000011110111;
20'b00011000110010011101: color_data = 12'b000011110111;
20'b00011000110010011110: color_data = 12'b000011110111;
20'b00011000110010011111: color_data = 12'b000011110111;
20'b00011000110010100001: color_data = 12'b000011110111;
20'b00011000110010100010: color_data = 12'b000011110111;
20'b00011000110010100011: color_data = 12'b000011110111;
20'b00011000110010100100: color_data = 12'b000011110111;
20'b00011000110010100101: color_data = 12'b000011110111;
20'b00011000110010100110: color_data = 12'b000011110111;
20'b00011000110010100111: color_data = 12'b000011110111;
20'b00011000110010101000: color_data = 12'b000011110111;
20'b00011000110010101001: color_data = 12'b000011110111;
20'b00011000110010101010: color_data = 12'b000011110111;
20'b00011000110100011010: color_data = 12'b000000001111;
20'b00011000110100011011: color_data = 12'b000000001111;
20'b00011000110100011100: color_data = 12'b000000001111;
20'b00011000110100011101: color_data = 12'b000000001111;
20'b00011000110100011110: color_data = 12'b000000001111;
20'b00011000110100011111: color_data = 12'b000000001111;
20'b00011000110100100000: color_data = 12'b000000001111;
20'b00011000110100100001: color_data = 12'b000000001111;
20'b00011000110100100010: color_data = 12'b000000001111;
20'b00011000110100100011: color_data = 12'b000000001111;
20'b00011000110110011110: color_data = 12'b000011110111;
20'b00011000110110011111: color_data = 12'b000011110111;
20'b00011000110110100000: color_data = 12'b000011110111;
20'b00011000110110100001: color_data = 12'b000011110111;
20'b00011000110110100010: color_data = 12'b000011110111;
20'b00011000110110100011: color_data = 12'b000011110111;
20'b00011000110110100100: color_data = 12'b000011110111;
20'b00011000110110100101: color_data = 12'b000011110111;
20'b00011000110110100110: color_data = 12'b000011110111;
20'b00011000110110100111: color_data = 12'b000011110111;
20'b00011001000010010110: color_data = 12'b000011110111;
20'b00011001000010010111: color_data = 12'b000011110111;
20'b00011001000010011000: color_data = 12'b000011110111;
20'b00011001000010011001: color_data = 12'b000011110111;
20'b00011001000010011010: color_data = 12'b000011110111;
20'b00011001000010011011: color_data = 12'b000011110111;
20'b00011001000010011100: color_data = 12'b000011110111;
20'b00011001000010011101: color_data = 12'b000011110111;
20'b00011001000010011110: color_data = 12'b000011110111;
20'b00011001000010011111: color_data = 12'b000011110111;
20'b00011001000010100001: color_data = 12'b000011110111;
20'b00011001000010100010: color_data = 12'b000011110111;
20'b00011001000010100011: color_data = 12'b000011110111;
20'b00011001000010100100: color_data = 12'b000011110111;
20'b00011001000010100101: color_data = 12'b000011110111;
20'b00011001000010100110: color_data = 12'b000011110111;
20'b00011001000010100111: color_data = 12'b000011110111;
20'b00011001000010101000: color_data = 12'b000011110111;
20'b00011001000010101001: color_data = 12'b000011110111;
20'b00011001000010101010: color_data = 12'b000011110111;
20'b00011001000100011010: color_data = 12'b000000001111;
20'b00011001000100011011: color_data = 12'b000000001111;
20'b00011001000100011100: color_data = 12'b000000001111;
20'b00011001000100011101: color_data = 12'b000000001111;
20'b00011001000100011110: color_data = 12'b000000001111;
20'b00011001000100011111: color_data = 12'b000000001111;
20'b00011001000100100000: color_data = 12'b000000001111;
20'b00011001000100100001: color_data = 12'b000000001111;
20'b00011001000100100010: color_data = 12'b000000001111;
20'b00011001000100100011: color_data = 12'b000000001111;
20'b00011001000110011110: color_data = 12'b000011110111;
20'b00011001000110011111: color_data = 12'b000011110111;
20'b00011001000110100000: color_data = 12'b000011110111;
20'b00011001000110100001: color_data = 12'b000011110111;
20'b00011001000110100010: color_data = 12'b000011110111;
20'b00011001000110100011: color_data = 12'b000011110111;
20'b00011001000110100100: color_data = 12'b000011110111;
20'b00011001000110100101: color_data = 12'b000011110111;
20'b00011001000110100110: color_data = 12'b000011110111;
20'b00011001000110100111: color_data = 12'b000011110111;
20'b00011001010010010110: color_data = 12'b000011110111;
20'b00011001010010010111: color_data = 12'b000011110111;
20'b00011001010010011000: color_data = 12'b000011110111;
20'b00011001010010011001: color_data = 12'b000011110111;
20'b00011001010010011010: color_data = 12'b000011110111;
20'b00011001010010011011: color_data = 12'b000011110111;
20'b00011001010010011100: color_data = 12'b000011110111;
20'b00011001010010011101: color_data = 12'b000011110111;
20'b00011001010010011110: color_data = 12'b000011110111;
20'b00011001010010011111: color_data = 12'b000011110111;
20'b00011001010010100001: color_data = 12'b000011110111;
20'b00011001010010100010: color_data = 12'b000011110111;
20'b00011001010010100011: color_data = 12'b000011110111;
20'b00011001010010100100: color_data = 12'b000011110111;
20'b00011001010010100101: color_data = 12'b000011110111;
20'b00011001010010100110: color_data = 12'b000011110111;
20'b00011001010010100111: color_data = 12'b000011110111;
20'b00011001010010101000: color_data = 12'b000011110111;
20'b00011001010010101001: color_data = 12'b000011110111;
20'b00011001010010101010: color_data = 12'b000011110111;
20'b00011001010100011010: color_data = 12'b000000001111;
20'b00011001010100011011: color_data = 12'b000000001111;
20'b00011001010100011100: color_data = 12'b000000001111;
20'b00011001010100011101: color_data = 12'b000000001111;
20'b00011001010100011110: color_data = 12'b000000001111;
20'b00011001010100011111: color_data = 12'b000000001111;
20'b00011001010100100000: color_data = 12'b000000001111;
20'b00011001010100100001: color_data = 12'b000000001111;
20'b00011001010100100010: color_data = 12'b000000001111;
20'b00011001010100100011: color_data = 12'b000000001111;
20'b00011001010110011110: color_data = 12'b000011110111;
20'b00011001010110011111: color_data = 12'b000011110111;
20'b00011001010110100000: color_data = 12'b000011110111;
20'b00011001010110100001: color_data = 12'b000011110111;
20'b00011001010110100010: color_data = 12'b000011110111;
20'b00011001010110100011: color_data = 12'b000011110111;
20'b00011001010110100100: color_data = 12'b000011110111;
20'b00011001010110100101: color_data = 12'b000011110111;
20'b00011001010110100110: color_data = 12'b000011110111;
20'b00011001010110100111: color_data = 12'b000011110111;
20'b00011001100010010110: color_data = 12'b000011110111;
20'b00011001100010010111: color_data = 12'b000011110111;
20'b00011001100010011000: color_data = 12'b000011110111;
20'b00011001100010011001: color_data = 12'b000011110111;
20'b00011001100010011010: color_data = 12'b000011110111;
20'b00011001100010011011: color_data = 12'b000011110111;
20'b00011001100010011100: color_data = 12'b000011110111;
20'b00011001100010011101: color_data = 12'b000011110111;
20'b00011001100010011110: color_data = 12'b000011110111;
20'b00011001100010011111: color_data = 12'b000011110111;
20'b00011001100010100001: color_data = 12'b000011110111;
20'b00011001100010100010: color_data = 12'b000011110111;
20'b00011001100010100011: color_data = 12'b000011110111;
20'b00011001100010100100: color_data = 12'b000011110111;
20'b00011001100010100101: color_data = 12'b000011110111;
20'b00011001100010100110: color_data = 12'b000011110111;
20'b00011001100010100111: color_data = 12'b000011110111;
20'b00011001100010101000: color_data = 12'b000011110111;
20'b00011001100010101001: color_data = 12'b000011110111;
20'b00011001100010101010: color_data = 12'b000011110111;
20'b00011001100100011010: color_data = 12'b000000001111;
20'b00011001100100011011: color_data = 12'b000000001111;
20'b00011001100100011100: color_data = 12'b000000001111;
20'b00011001100100011101: color_data = 12'b000000001111;
20'b00011001100100011110: color_data = 12'b000000001111;
20'b00011001100100011111: color_data = 12'b000000001111;
20'b00011001100100100000: color_data = 12'b000000001111;
20'b00011001100100100001: color_data = 12'b000000001111;
20'b00011001100100100010: color_data = 12'b000000001111;
20'b00011001100100100011: color_data = 12'b000000001111;
20'b00011001100110011110: color_data = 12'b000011110111;
20'b00011001100110011111: color_data = 12'b000011110111;
20'b00011001100110100000: color_data = 12'b000011110111;
20'b00011001100110100001: color_data = 12'b000011110111;
20'b00011001100110100010: color_data = 12'b000011110111;
20'b00011001100110100011: color_data = 12'b000011110111;
20'b00011001100110100100: color_data = 12'b000011110111;
20'b00011001100110100101: color_data = 12'b000011110111;
20'b00011001100110100110: color_data = 12'b000011110111;
20'b00011001100110100111: color_data = 12'b000011110111;
20'b00011001110110011110: color_data = 12'b000011110111;
20'b00011001110110011111: color_data = 12'b000011110111;
20'b00011001110110100000: color_data = 12'b000011110111;
20'b00011001110110100001: color_data = 12'b000011110111;
20'b00011001110110100010: color_data = 12'b000011110111;
20'b00011001110110100011: color_data = 12'b000011110111;
20'b00011001110110100100: color_data = 12'b000011110111;
20'b00011001110110100101: color_data = 12'b000011110111;
20'b00011001110110100110: color_data = 12'b000011110111;
20'b00011001110110100111: color_data = 12'b000011110111;
20'b00011010000101000110: color_data = 12'b111100000000;
20'b00011010000101000111: color_data = 12'b111100000000;
20'b00011010000101001000: color_data = 12'b111100000000;
20'b00011010000101001001: color_data = 12'b111100000000;
20'b00011010000101001010: color_data = 12'b111100000000;
20'b00011010000101001011: color_data = 12'b111100000000;
20'b00011010000101001100: color_data = 12'b111100000000;
20'b00011010000101001101: color_data = 12'b111100000000;
20'b00011010000101001110: color_data = 12'b111100000000;
20'b00011010000101001111: color_data = 12'b111100000000;
20'b00011010000101010001: color_data = 12'b111100000000;
20'b00011010000101010010: color_data = 12'b111100000000;
20'b00011010000101010011: color_data = 12'b111100000000;
20'b00011010000101010100: color_data = 12'b111100000000;
20'b00011010000101010101: color_data = 12'b111100000000;
20'b00011010000101010110: color_data = 12'b111100000000;
20'b00011010000101010111: color_data = 12'b111100000000;
20'b00011010000101011000: color_data = 12'b111100000000;
20'b00011010000101011001: color_data = 12'b111100000000;
20'b00011010000101011010: color_data = 12'b111100000000;
20'b00011010000110011110: color_data = 12'b000011110111;
20'b00011010000110011111: color_data = 12'b000011110111;
20'b00011010000110100000: color_data = 12'b000011110111;
20'b00011010000110100001: color_data = 12'b000011110111;
20'b00011010000110100010: color_data = 12'b000011110111;
20'b00011010000110100011: color_data = 12'b000011110111;
20'b00011010000110100100: color_data = 12'b000011110111;
20'b00011010000110100101: color_data = 12'b000011110111;
20'b00011010000110100110: color_data = 12'b000011110111;
20'b00011010000110100111: color_data = 12'b000011110111;
20'b00011010010101000110: color_data = 12'b111100000000;
20'b00011010010101000111: color_data = 12'b111100000000;
20'b00011010010101001000: color_data = 12'b111100000000;
20'b00011010010101001001: color_data = 12'b111100000000;
20'b00011010010101001010: color_data = 12'b111100000000;
20'b00011010010101001011: color_data = 12'b111100000000;
20'b00011010010101001100: color_data = 12'b111100000000;
20'b00011010010101001101: color_data = 12'b111100000000;
20'b00011010010101001110: color_data = 12'b111100000000;
20'b00011010010101001111: color_data = 12'b111100000000;
20'b00011010010101010001: color_data = 12'b111100000000;
20'b00011010010101010010: color_data = 12'b111100000000;
20'b00011010010101010011: color_data = 12'b111100000000;
20'b00011010010101010100: color_data = 12'b111100000000;
20'b00011010010101010101: color_data = 12'b111100000000;
20'b00011010010101010110: color_data = 12'b111100000000;
20'b00011010010101010111: color_data = 12'b111100000000;
20'b00011010010101011000: color_data = 12'b111100000000;
20'b00011010010101011001: color_data = 12'b111100000000;
20'b00011010010101011010: color_data = 12'b111100000000;
20'b00011010010110011110: color_data = 12'b000011110111;
20'b00011010010110011111: color_data = 12'b000011110111;
20'b00011010010110100000: color_data = 12'b000011110111;
20'b00011010010110100001: color_data = 12'b000011110111;
20'b00011010010110100010: color_data = 12'b000011110111;
20'b00011010010110100011: color_data = 12'b000011110111;
20'b00011010010110100100: color_data = 12'b000011110111;
20'b00011010010110100101: color_data = 12'b000011110111;
20'b00011010010110100110: color_data = 12'b000011110111;
20'b00011010010110100111: color_data = 12'b000011110111;
20'b00011010100101000110: color_data = 12'b111100000000;
20'b00011010100101000111: color_data = 12'b111100000000;
20'b00011010100101001000: color_data = 12'b111100000000;
20'b00011010100101001001: color_data = 12'b111100000000;
20'b00011010100101001010: color_data = 12'b111100000000;
20'b00011010100101001011: color_data = 12'b111100000000;
20'b00011010100101001100: color_data = 12'b111100000000;
20'b00011010100101001101: color_data = 12'b111100000000;
20'b00011010100101001110: color_data = 12'b111100000000;
20'b00011010100101001111: color_data = 12'b111100000000;
20'b00011010100101010001: color_data = 12'b111100000000;
20'b00011010100101010010: color_data = 12'b111100000000;
20'b00011010100101010011: color_data = 12'b111100000000;
20'b00011010100101010100: color_data = 12'b111100000000;
20'b00011010100101010101: color_data = 12'b111100000000;
20'b00011010100101010110: color_data = 12'b111100000000;
20'b00011010100101010111: color_data = 12'b111100000000;
20'b00011010100101011000: color_data = 12'b111100000000;
20'b00011010100101011001: color_data = 12'b111100000000;
20'b00011010100101011010: color_data = 12'b111100000000;
20'b00011010110101000110: color_data = 12'b111100000000;
20'b00011010110101000111: color_data = 12'b111100000000;
20'b00011010110101001000: color_data = 12'b111100000000;
20'b00011010110101001001: color_data = 12'b111100000000;
20'b00011010110101001010: color_data = 12'b111100000000;
20'b00011010110101001011: color_data = 12'b111100000000;
20'b00011010110101001100: color_data = 12'b111100000000;
20'b00011010110101001101: color_data = 12'b111100000000;
20'b00011010110101001110: color_data = 12'b111100000000;
20'b00011010110101001111: color_data = 12'b111100000000;
20'b00011010110101010001: color_data = 12'b111100000000;
20'b00011010110101010010: color_data = 12'b111100000000;
20'b00011010110101010011: color_data = 12'b111100000000;
20'b00011010110101010100: color_data = 12'b111100000000;
20'b00011010110101010101: color_data = 12'b111100000000;
20'b00011010110101010110: color_data = 12'b111100000000;
20'b00011010110101010111: color_data = 12'b111100000000;
20'b00011010110101011000: color_data = 12'b111100000000;
20'b00011010110101011001: color_data = 12'b111100000000;
20'b00011010110101011010: color_data = 12'b111100000000;
20'b00011010110110011110: color_data = 12'b000011110111;
20'b00011010110110011111: color_data = 12'b000011110111;
20'b00011010110110100000: color_data = 12'b000011110111;
20'b00011010110110100001: color_data = 12'b000011110111;
20'b00011010110110100010: color_data = 12'b000011110111;
20'b00011010110110100011: color_data = 12'b000011110111;
20'b00011010110110100100: color_data = 12'b000011110111;
20'b00011010110110100101: color_data = 12'b000011110111;
20'b00011010110110100110: color_data = 12'b000011110111;
20'b00011010110110100111: color_data = 12'b000011110111;
20'b00011011000101000110: color_data = 12'b111100000000;
20'b00011011000101000111: color_data = 12'b111100000000;
20'b00011011000101001000: color_data = 12'b111100000000;
20'b00011011000101001001: color_data = 12'b111100000000;
20'b00011011000101001010: color_data = 12'b111100000000;
20'b00011011000101001011: color_data = 12'b111100000000;
20'b00011011000101001100: color_data = 12'b111100000000;
20'b00011011000101001101: color_data = 12'b111100000000;
20'b00011011000101001110: color_data = 12'b111100000000;
20'b00011011000101001111: color_data = 12'b111100000000;
20'b00011011000101010001: color_data = 12'b111100000000;
20'b00011011000101010010: color_data = 12'b111100000000;
20'b00011011000101010011: color_data = 12'b111100000000;
20'b00011011000101010100: color_data = 12'b111100000000;
20'b00011011000101010101: color_data = 12'b111100000000;
20'b00011011000101010110: color_data = 12'b111100000000;
20'b00011011000101010111: color_data = 12'b111100000000;
20'b00011011000101011000: color_data = 12'b111100000000;
20'b00011011000101011001: color_data = 12'b111100000000;
20'b00011011000101011010: color_data = 12'b111100000000;
20'b00011011000110011110: color_data = 12'b000011110111;
20'b00011011000110011111: color_data = 12'b000011110111;
20'b00011011000110100000: color_data = 12'b000011110111;
20'b00011011000110100001: color_data = 12'b000011110111;
20'b00011011000110100010: color_data = 12'b000011110111;
20'b00011011000110100011: color_data = 12'b000011110111;
20'b00011011000110100100: color_data = 12'b000011110111;
20'b00011011000110100101: color_data = 12'b000011110111;
20'b00011011000110100110: color_data = 12'b000011110111;
20'b00011011000110100111: color_data = 12'b000011110111;
20'b00011011010101000110: color_data = 12'b111100000000;
20'b00011011010101000111: color_data = 12'b111100000000;
20'b00011011010101001000: color_data = 12'b111100000000;
20'b00011011010101001001: color_data = 12'b111100000000;
20'b00011011010101001010: color_data = 12'b111100000000;
20'b00011011010101001011: color_data = 12'b111100000000;
20'b00011011010101001100: color_data = 12'b111100000000;
20'b00011011010101001101: color_data = 12'b111100000000;
20'b00011011010101001110: color_data = 12'b111100000000;
20'b00011011010101001111: color_data = 12'b111100000000;
20'b00011011010101010001: color_data = 12'b111100000000;
20'b00011011010101010010: color_data = 12'b111100000000;
20'b00011011010101010011: color_data = 12'b111100000000;
20'b00011011010101010100: color_data = 12'b111100000000;
20'b00011011010101010101: color_data = 12'b111100000000;
20'b00011011010101010110: color_data = 12'b111100000000;
20'b00011011010101010111: color_data = 12'b111100000000;
20'b00011011010101011000: color_data = 12'b111100000000;
20'b00011011010101011001: color_data = 12'b111100000000;
20'b00011011010101011010: color_data = 12'b111100000000;
20'b00011011010110011110: color_data = 12'b000011110111;
20'b00011011010110011111: color_data = 12'b000011110111;
20'b00011011010110100000: color_data = 12'b000011110111;
20'b00011011010110100001: color_data = 12'b000011110111;
20'b00011011010110100010: color_data = 12'b000011110111;
20'b00011011010110100011: color_data = 12'b000011110111;
20'b00011011010110100100: color_data = 12'b000011110111;
20'b00011011010110100101: color_data = 12'b000011110111;
20'b00011011010110100110: color_data = 12'b000011110111;
20'b00011011010110100111: color_data = 12'b000011110111;
20'b00011011100101000110: color_data = 12'b111100000000;
20'b00011011100101000111: color_data = 12'b111100000000;
20'b00011011100101001000: color_data = 12'b111100000000;
20'b00011011100101001001: color_data = 12'b111100000000;
20'b00011011100101001010: color_data = 12'b111100000000;
20'b00011011100101001011: color_data = 12'b111100000000;
20'b00011011100101001100: color_data = 12'b111100000000;
20'b00011011100101001101: color_data = 12'b111100000000;
20'b00011011100101001110: color_data = 12'b111100000000;
20'b00011011100101001111: color_data = 12'b111100000000;
20'b00011011100101010001: color_data = 12'b111100000000;
20'b00011011100101010010: color_data = 12'b111100000000;
20'b00011011100101010011: color_data = 12'b111100000000;
20'b00011011100101010100: color_data = 12'b111100000000;
20'b00011011100101010101: color_data = 12'b111100000000;
20'b00011011100101010110: color_data = 12'b111100000000;
20'b00011011100101010111: color_data = 12'b111100000000;
20'b00011011100101011000: color_data = 12'b111100000000;
20'b00011011100101011001: color_data = 12'b111100000000;
20'b00011011100101011010: color_data = 12'b111100000000;
20'b00011011100110011110: color_data = 12'b000011110111;
20'b00011011100110011111: color_data = 12'b000011110111;
20'b00011011100110100000: color_data = 12'b000011110111;
20'b00011011100110100001: color_data = 12'b000011110111;
20'b00011011100110100010: color_data = 12'b000011110111;
20'b00011011100110100011: color_data = 12'b000011110111;
20'b00011011100110100100: color_data = 12'b000011110111;
20'b00011011100110100101: color_data = 12'b000011110111;
20'b00011011100110100110: color_data = 12'b000011110111;
20'b00011011100110100111: color_data = 12'b000011110111;
20'b00011011110101000110: color_data = 12'b111100000000;
20'b00011011110101000111: color_data = 12'b111100000000;
20'b00011011110101001000: color_data = 12'b111100000000;
20'b00011011110101001001: color_data = 12'b111100000000;
20'b00011011110101001010: color_data = 12'b111100000000;
20'b00011011110101001011: color_data = 12'b111100000000;
20'b00011011110101001100: color_data = 12'b111100000000;
20'b00011011110101001101: color_data = 12'b111100000000;
20'b00011011110101001110: color_data = 12'b111100000000;
20'b00011011110101001111: color_data = 12'b111100000000;
20'b00011011110101010001: color_data = 12'b111100000000;
20'b00011011110101010010: color_data = 12'b111100000000;
20'b00011011110101010011: color_data = 12'b111100000000;
20'b00011011110101010100: color_data = 12'b111100000000;
20'b00011011110101010101: color_data = 12'b111100000000;
20'b00011011110101010110: color_data = 12'b111100000000;
20'b00011011110101010111: color_data = 12'b111100000000;
20'b00011011110101011000: color_data = 12'b111100000000;
20'b00011011110101011001: color_data = 12'b111100000000;
20'b00011011110101011010: color_data = 12'b111100000000;
20'b00011011110110011110: color_data = 12'b000011110111;
20'b00011011110110011111: color_data = 12'b000011110111;
20'b00011011110110100000: color_data = 12'b000011110111;
20'b00011011110110100001: color_data = 12'b000011110111;
20'b00011011110110100010: color_data = 12'b000011110111;
20'b00011011110110100011: color_data = 12'b000011110111;
20'b00011011110110100100: color_data = 12'b000011110111;
20'b00011011110110100101: color_data = 12'b000011110111;
20'b00011011110110100110: color_data = 12'b000011110111;
20'b00011011110110100111: color_data = 12'b000011110111;
20'b00011100000101000110: color_data = 12'b111100000000;
20'b00011100000101000111: color_data = 12'b111100000000;
20'b00011100000101001000: color_data = 12'b111100000000;
20'b00011100000101001001: color_data = 12'b111100000000;
20'b00011100000101001010: color_data = 12'b111100000000;
20'b00011100000101001011: color_data = 12'b111100000000;
20'b00011100000101001100: color_data = 12'b111100000000;
20'b00011100000101001101: color_data = 12'b111100000000;
20'b00011100000101001110: color_data = 12'b111100000000;
20'b00011100000101001111: color_data = 12'b111100000000;
20'b00011100000101010001: color_data = 12'b111100000000;
20'b00011100000101010010: color_data = 12'b111100000000;
20'b00011100000101010011: color_data = 12'b111100000000;
20'b00011100000101010100: color_data = 12'b111100000000;
20'b00011100000101010101: color_data = 12'b111100000000;
20'b00011100000101010110: color_data = 12'b111100000000;
20'b00011100000101010111: color_data = 12'b111100000000;
20'b00011100000101011000: color_data = 12'b111100000000;
20'b00011100000101011001: color_data = 12'b111100000000;
20'b00011100000101011010: color_data = 12'b111100000000;
20'b00011100000110011110: color_data = 12'b000011110111;
20'b00011100000110011111: color_data = 12'b000011110111;
20'b00011100000110100000: color_data = 12'b000011110111;
20'b00011100000110100001: color_data = 12'b000011110111;
20'b00011100000110100010: color_data = 12'b000011110111;
20'b00011100000110100011: color_data = 12'b000011110111;
20'b00011100000110100100: color_data = 12'b000011110111;
20'b00011100000110100101: color_data = 12'b000011110111;
20'b00011100000110100110: color_data = 12'b000011110111;
20'b00011100000110100111: color_data = 12'b000011110111;
20'b00011100010101000110: color_data = 12'b111100000000;
20'b00011100010101000111: color_data = 12'b111100000000;
20'b00011100010101001000: color_data = 12'b111100000000;
20'b00011100010101001001: color_data = 12'b111100000000;
20'b00011100010101001010: color_data = 12'b111100000000;
20'b00011100010101001011: color_data = 12'b111100000000;
20'b00011100010101001100: color_data = 12'b111100000000;
20'b00011100010101001101: color_data = 12'b111100000000;
20'b00011100010101001110: color_data = 12'b111100000000;
20'b00011100010101001111: color_data = 12'b111100000000;
20'b00011100010101010001: color_data = 12'b111100000000;
20'b00011100010101010010: color_data = 12'b111100000000;
20'b00011100010101010011: color_data = 12'b111100000000;
20'b00011100010101010100: color_data = 12'b111100000000;
20'b00011100010101010101: color_data = 12'b111100000000;
20'b00011100010101010110: color_data = 12'b111100000000;
20'b00011100010101010111: color_data = 12'b111100000000;
20'b00011100010101011000: color_data = 12'b111100000000;
20'b00011100010101011001: color_data = 12'b111100000000;
20'b00011100010101011010: color_data = 12'b111100000000;
20'b00011100010110011110: color_data = 12'b000011110111;
20'b00011100010110011111: color_data = 12'b000011110111;
20'b00011100010110100000: color_data = 12'b000011110111;
20'b00011100010110100001: color_data = 12'b000011110111;
20'b00011100010110100010: color_data = 12'b000011110111;
20'b00011100010110100011: color_data = 12'b000011110111;
20'b00011100010110100100: color_data = 12'b000011110111;
20'b00011100010110100101: color_data = 12'b000011110111;
20'b00011100010110100110: color_data = 12'b000011110111;
20'b00011100010110100111: color_data = 12'b000011110111;
20'b00011100100110011110: color_data = 12'b000011110111;
20'b00011100100110011111: color_data = 12'b000011110111;
20'b00011100100110100000: color_data = 12'b000011110111;
20'b00011100100110100001: color_data = 12'b000011110111;
20'b00011100100110100010: color_data = 12'b000011110111;
20'b00011100100110100011: color_data = 12'b000011110111;
20'b00011100100110100100: color_data = 12'b000011110111;
20'b00011100100110100101: color_data = 12'b000011110111;
20'b00011100100110100110: color_data = 12'b000011110111;
20'b00011100100110100111: color_data = 12'b000011110111;
20'b00011100110010101100: color_data = 12'b111011101110;
20'b00011100110010101101: color_data = 12'b111011101110;
20'b00011100110010101110: color_data = 12'b111011101110;
20'b00011100110010101111: color_data = 12'b111011101110;
20'b00011100110010110000: color_data = 12'b111011101110;
20'b00011100110010110001: color_data = 12'b111011101110;
20'b00011100110010110010: color_data = 12'b111011101110;
20'b00011100110010110011: color_data = 12'b111011101110;
20'b00011100110010110100: color_data = 12'b111011101110;
20'b00011100110010110101: color_data = 12'b111011101110;
20'b00011100110010110111: color_data = 12'b111011101110;
20'b00011100110010111000: color_data = 12'b111011101110;
20'b00011100110010111001: color_data = 12'b111011101110;
20'b00011100110010111010: color_data = 12'b111011101110;
20'b00011100110010111011: color_data = 12'b111011101110;
20'b00011100110010111100: color_data = 12'b111011101110;
20'b00011100110010111101: color_data = 12'b111011101110;
20'b00011100110010111110: color_data = 12'b111011101110;
20'b00011100110010111111: color_data = 12'b111011101110;
20'b00011100110011000000: color_data = 12'b111011101110;
20'b00011100110011000010: color_data = 12'b111011101110;
20'b00011100110011000011: color_data = 12'b111011101110;
20'b00011100110011000100: color_data = 12'b111011101110;
20'b00011100110011000101: color_data = 12'b111011101110;
20'b00011100110011000110: color_data = 12'b111011101110;
20'b00011100110011000111: color_data = 12'b111011101110;
20'b00011100110011001000: color_data = 12'b111011101110;
20'b00011100110011001001: color_data = 12'b111011101110;
20'b00011100110011001010: color_data = 12'b111011101110;
20'b00011100110011001011: color_data = 12'b111011101110;
20'b00011100110011001101: color_data = 12'b111011101110;
20'b00011100110011001110: color_data = 12'b111011101110;
20'b00011100110011001111: color_data = 12'b111011101110;
20'b00011100110011010000: color_data = 12'b111011101110;
20'b00011100110011010001: color_data = 12'b111011101110;
20'b00011100110011010010: color_data = 12'b111011101110;
20'b00011100110011010011: color_data = 12'b111011101110;
20'b00011100110011010100: color_data = 12'b111011101110;
20'b00011100110011010101: color_data = 12'b111011101110;
20'b00011100110011010110: color_data = 12'b111011101110;
20'b00011100110100000100: color_data = 12'b111011101110;
20'b00011100110100000101: color_data = 12'b111011101110;
20'b00011100110100000110: color_data = 12'b111011101110;
20'b00011100110100000111: color_data = 12'b111011101110;
20'b00011100110100001000: color_data = 12'b111011101110;
20'b00011100110100001001: color_data = 12'b111011101110;
20'b00011100110100001010: color_data = 12'b111011101110;
20'b00011100110100001011: color_data = 12'b111011101110;
20'b00011100110100001100: color_data = 12'b111011101110;
20'b00011100110100001101: color_data = 12'b111011101110;
20'b00011100110101010001: color_data = 12'b111100000000;
20'b00011100110101010010: color_data = 12'b111100000000;
20'b00011100110101010011: color_data = 12'b111100000000;
20'b00011100110101010100: color_data = 12'b111100000000;
20'b00011100110101010101: color_data = 12'b111100000000;
20'b00011100110101010110: color_data = 12'b111100000000;
20'b00011100110101010111: color_data = 12'b111100000000;
20'b00011100110101011000: color_data = 12'b111100000000;
20'b00011100110101011001: color_data = 12'b111100000000;
20'b00011100110101011010: color_data = 12'b111100000000;
20'b00011100110101011100: color_data = 12'b111100000000;
20'b00011100110101011101: color_data = 12'b111100000000;
20'b00011100110101011110: color_data = 12'b111100000000;
20'b00011100110101011111: color_data = 12'b111100000000;
20'b00011100110101100000: color_data = 12'b111100000000;
20'b00011100110101100001: color_data = 12'b111100000000;
20'b00011100110101100010: color_data = 12'b111100000000;
20'b00011100110101100011: color_data = 12'b111100000000;
20'b00011100110101100100: color_data = 12'b111100000000;
20'b00011100110101100101: color_data = 12'b111100000000;
20'b00011100110101111101: color_data = 12'b111011101110;
20'b00011100110101111110: color_data = 12'b111011101110;
20'b00011100110101111111: color_data = 12'b111011101110;
20'b00011100110110000000: color_data = 12'b111011101110;
20'b00011100110110000001: color_data = 12'b111011101110;
20'b00011100110110000010: color_data = 12'b111011101110;
20'b00011100110110000011: color_data = 12'b111011101110;
20'b00011100110110000100: color_data = 12'b111011101110;
20'b00011100110110000101: color_data = 12'b111011101110;
20'b00011100110110000110: color_data = 12'b111011101110;
20'b00011100110110001000: color_data = 12'b111011101110;
20'b00011100110110001001: color_data = 12'b111011101110;
20'b00011100110110001010: color_data = 12'b111011101110;
20'b00011100110110001011: color_data = 12'b111011101110;
20'b00011100110110001100: color_data = 12'b111011101110;
20'b00011100110110001101: color_data = 12'b111011101110;
20'b00011100110110001110: color_data = 12'b111011101110;
20'b00011100110110001111: color_data = 12'b111011101110;
20'b00011100110110010000: color_data = 12'b111011101110;
20'b00011100110110010001: color_data = 12'b111011101110;
20'b00011100110110011110: color_data = 12'b000011110111;
20'b00011100110110011111: color_data = 12'b000011110111;
20'b00011100110110100000: color_data = 12'b000011110111;
20'b00011100110110100001: color_data = 12'b000011110111;
20'b00011100110110100010: color_data = 12'b000011110111;
20'b00011100110110100011: color_data = 12'b000011110111;
20'b00011100110110100100: color_data = 12'b000011110111;
20'b00011100110110100101: color_data = 12'b000011110111;
20'b00011100110110100110: color_data = 12'b000011110111;
20'b00011100110110100111: color_data = 12'b000011110111;
20'b00011101000010101100: color_data = 12'b111011101110;
20'b00011101000010101101: color_data = 12'b111011101110;
20'b00011101000010101110: color_data = 12'b111011101110;
20'b00011101000010101111: color_data = 12'b111011101110;
20'b00011101000010110000: color_data = 12'b111011101110;
20'b00011101000010110001: color_data = 12'b111011101110;
20'b00011101000010110010: color_data = 12'b111011101110;
20'b00011101000010110011: color_data = 12'b111011101110;
20'b00011101000010110100: color_data = 12'b111011101110;
20'b00011101000010110101: color_data = 12'b111011101110;
20'b00011101000010110111: color_data = 12'b111011101110;
20'b00011101000010111000: color_data = 12'b111011101110;
20'b00011101000010111001: color_data = 12'b111011101110;
20'b00011101000010111010: color_data = 12'b111011101110;
20'b00011101000010111011: color_data = 12'b111011101110;
20'b00011101000010111100: color_data = 12'b111011101110;
20'b00011101000010111101: color_data = 12'b111011101110;
20'b00011101000010111110: color_data = 12'b111011101110;
20'b00011101000010111111: color_data = 12'b111011101110;
20'b00011101000011000000: color_data = 12'b111011101110;
20'b00011101000011000010: color_data = 12'b111011101110;
20'b00011101000011000011: color_data = 12'b111011101110;
20'b00011101000011000100: color_data = 12'b111011101110;
20'b00011101000011000101: color_data = 12'b111011101110;
20'b00011101000011000110: color_data = 12'b111011101110;
20'b00011101000011000111: color_data = 12'b111011101110;
20'b00011101000011001000: color_data = 12'b111011101110;
20'b00011101000011001001: color_data = 12'b111011101110;
20'b00011101000011001010: color_data = 12'b111011101110;
20'b00011101000011001011: color_data = 12'b111011101110;
20'b00011101000011001101: color_data = 12'b111011101110;
20'b00011101000011001110: color_data = 12'b111011101110;
20'b00011101000011001111: color_data = 12'b111011101110;
20'b00011101000011010000: color_data = 12'b111011101110;
20'b00011101000011010001: color_data = 12'b111011101110;
20'b00011101000011010010: color_data = 12'b111011101110;
20'b00011101000011010011: color_data = 12'b111011101110;
20'b00011101000011010100: color_data = 12'b111011101110;
20'b00011101000011010101: color_data = 12'b111011101110;
20'b00011101000011010110: color_data = 12'b111011101110;
20'b00011101000100000100: color_data = 12'b111011101110;
20'b00011101000100000101: color_data = 12'b111011101110;
20'b00011101000100000110: color_data = 12'b111011101110;
20'b00011101000100000111: color_data = 12'b111011101110;
20'b00011101000100001000: color_data = 12'b111011101110;
20'b00011101000100001001: color_data = 12'b111011101110;
20'b00011101000100001010: color_data = 12'b111011101110;
20'b00011101000100001011: color_data = 12'b111011101110;
20'b00011101000100001100: color_data = 12'b111011101110;
20'b00011101000100001101: color_data = 12'b111011101110;
20'b00011101000101010001: color_data = 12'b111100000000;
20'b00011101000101010010: color_data = 12'b111100000000;
20'b00011101000101010011: color_data = 12'b111100000000;
20'b00011101000101010100: color_data = 12'b111100000000;
20'b00011101000101010101: color_data = 12'b111100000000;
20'b00011101000101010110: color_data = 12'b111100000000;
20'b00011101000101010111: color_data = 12'b111100000000;
20'b00011101000101011000: color_data = 12'b111100000000;
20'b00011101000101011001: color_data = 12'b111100000000;
20'b00011101000101011010: color_data = 12'b111100000000;
20'b00011101000101011100: color_data = 12'b111100000000;
20'b00011101000101011101: color_data = 12'b111100000000;
20'b00011101000101011110: color_data = 12'b111100000000;
20'b00011101000101011111: color_data = 12'b111100000000;
20'b00011101000101100000: color_data = 12'b111100000000;
20'b00011101000101100001: color_data = 12'b111100000000;
20'b00011101000101100010: color_data = 12'b111100000000;
20'b00011101000101100011: color_data = 12'b111100000000;
20'b00011101000101100100: color_data = 12'b111100000000;
20'b00011101000101100101: color_data = 12'b111100000000;
20'b00011101000101111101: color_data = 12'b111011101110;
20'b00011101000101111110: color_data = 12'b111011101110;
20'b00011101000101111111: color_data = 12'b111011101110;
20'b00011101000110000000: color_data = 12'b111011101110;
20'b00011101000110000001: color_data = 12'b111011101110;
20'b00011101000110000010: color_data = 12'b111011101110;
20'b00011101000110000011: color_data = 12'b111011101110;
20'b00011101000110000100: color_data = 12'b111011101110;
20'b00011101000110000101: color_data = 12'b111011101110;
20'b00011101000110000110: color_data = 12'b111011101110;
20'b00011101000110001000: color_data = 12'b111011101110;
20'b00011101000110001001: color_data = 12'b111011101110;
20'b00011101000110001010: color_data = 12'b111011101110;
20'b00011101000110001011: color_data = 12'b111011101110;
20'b00011101000110001100: color_data = 12'b111011101110;
20'b00011101000110001101: color_data = 12'b111011101110;
20'b00011101000110001110: color_data = 12'b111011101110;
20'b00011101000110001111: color_data = 12'b111011101110;
20'b00011101000110010000: color_data = 12'b111011101110;
20'b00011101000110010001: color_data = 12'b111011101110;
20'b00011101010010101100: color_data = 12'b111011101110;
20'b00011101010010101101: color_data = 12'b111011101110;
20'b00011101010010101110: color_data = 12'b111011101110;
20'b00011101010010101111: color_data = 12'b111011101110;
20'b00011101010010110000: color_data = 12'b111011101110;
20'b00011101010010110001: color_data = 12'b111011101110;
20'b00011101010010110010: color_data = 12'b111011101110;
20'b00011101010010110011: color_data = 12'b111011101110;
20'b00011101010010110100: color_data = 12'b111011101110;
20'b00011101010010110101: color_data = 12'b111011101110;
20'b00011101010010110111: color_data = 12'b111011101110;
20'b00011101010010111000: color_data = 12'b111011101110;
20'b00011101010010111001: color_data = 12'b111011101110;
20'b00011101010010111010: color_data = 12'b111011101110;
20'b00011101010010111011: color_data = 12'b111011101110;
20'b00011101010010111100: color_data = 12'b111011101110;
20'b00011101010010111101: color_data = 12'b111011101110;
20'b00011101010010111110: color_data = 12'b111011101110;
20'b00011101010010111111: color_data = 12'b111011101110;
20'b00011101010011000000: color_data = 12'b111011101110;
20'b00011101010011000010: color_data = 12'b111011101110;
20'b00011101010011000011: color_data = 12'b111011101110;
20'b00011101010011000100: color_data = 12'b111011101110;
20'b00011101010011000101: color_data = 12'b111011101110;
20'b00011101010011000110: color_data = 12'b111011101110;
20'b00011101010011000111: color_data = 12'b111011101110;
20'b00011101010011001000: color_data = 12'b111011101110;
20'b00011101010011001001: color_data = 12'b111011101110;
20'b00011101010011001010: color_data = 12'b111011101110;
20'b00011101010011001011: color_data = 12'b111011101110;
20'b00011101010011001101: color_data = 12'b111011101110;
20'b00011101010011001110: color_data = 12'b111011101110;
20'b00011101010011001111: color_data = 12'b111011101110;
20'b00011101010011010000: color_data = 12'b111011101110;
20'b00011101010011010001: color_data = 12'b111011101110;
20'b00011101010011010010: color_data = 12'b111011101110;
20'b00011101010011010011: color_data = 12'b111011101110;
20'b00011101010011010100: color_data = 12'b111011101110;
20'b00011101010011010101: color_data = 12'b111011101110;
20'b00011101010011010110: color_data = 12'b111011101110;
20'b00011101010100000100: color_data = 12'b111011101110;
20'b00011101010100000101: color_data = 12'b111011101110;
20'b00011101010100000110: color_data = 12'b111011101110;
20'b00011101010100000111: color_data = 12'b111011101110;
20'b00011101010100001000: color_data = 12'b111011101110;
20'b00011101010100001001: color_data = 12'b111011101110;
20'b00011101010100001010: color_data = 12'b111011101110;
20'b00011101010100001011: color_data = 12'b111011101110;
20'b00011101010100001100: color_data = 12'b111011101110;
20'b00011101010100001101: color_data = 12'b111011101110;
20'b00011101010101010001: color_data = 12'b111100000000;
20'b00011101010101010010: color_data = 12'b111100000000;
20'b00011101010101010011: color_data = 12'b111100000000;
20'b00011101010101010100: color_data = 12'b111100000000;
20'b00011101010101010101: color_data = 12'b111100000000;
20'b00011101010101010110: color_data = 12'b111100000000;
20'b00011101010101010111: color_data = 12'b111100000000;
20'b00011101010101011000: color_data = 12'b111100000000;
20'b00011101010101011001: color_data = 12'b111100000000;
20'b00011101010101011010: color_data = 12'b111100000000;
20'b00011101010101011100: color_data = 12'b111100000000;
20'b00011101010101011101: color_data = 12'b111100000000;
20'b00011101010101011110: color_data = 12'b111100000000;
20'b00011101010101011111: color_data = 12'b111100000000;
20'b00011101010101100000: color_data = 12'b111100000000;
20'b00011101010101100001: color_data = 12'b111100000000;
20'b00011101010101100010: color_data = 12'b111100000000;
20'b00011101010101100011: color_data = 12'b111100000000;
20'b00011101010101100100: color_data = 12'b111100000000;
20'b00011101010101100101: color_data = 12'b111100000000;
20'b00011101010101111101: color_data = 12'b111011101110;
20'b00011101010101111110: color_data = 12'b111011101110;
20'b00011101010101111111: color_data = 12'b111011101110;
20'b00011101010110000000: color_data = 12'b111011101110;
20'b00011101010110000001: color_data = 12'b111011101110;
20'b00011101010110000010: color_data = 12'b111011101110;
20'b00011101010110000011: color_data = 12'b111011101110;
20'b00011101010110000100: color_data = 12'b111011101110;
20'b00011101010110000101: color_data = 12'b111011101110;
20'b00011101010110000110: color_data = 12'b111011101110;
20'b00011101010110001000: color_data = 12'b111011101110;
20'b00011101010110001001: color_data = 12'b111011101110;
20'b00011101010110001010: color_data = 12'b111011101110;
20'b00011101010110001011: color_data = 12'b111011101110;
20'b00011101010110001100: color_data = 12'b111011101110;
20'b00011101010110001101: color_data = 12'b111011101110;
20'b00011101010110001110: color_data = 12'b111011101110;
20'b00011101010110001111: color_data = 12'b111011101110;
20'b00011101010110010000: color_data = 12'b111011101110;
20'b00011101010110010001: color_data = 12'b111011101110;
20'b00011101010110110100: color_data = 12'b111011101110;
20'b00011101010110110101: color_data = 12'b111011101110;
20'b00011101010110110110: color_data = 12'b111011101110;
20'b00011101010110110111: color_data = 12'b111011101110;
20'b00011101010110111000: color_data = 12'b111011101110;
20'b00011101010110111001: color_data = 12'b111011101110;
20'b00011101010110111010: color_data = 12'b111011101110;
20'b00011101010110111011: color_data = 12'b111011101110;
20'b00011101010110111100: color_data = 12'b111011101110;
20'b00011101010110111101: color_data = 12'b111011101110;
20'b00011101010110111111: color_data = 12'b111011101110;
20'b00011101010111000000: color_data = 12'b111011101110;
20'b00011101010111000001: color_data = 12'b111011101110;
20'b00011101010111000010: color_data = 12'b111011101110;
20'b00011101010111000011: color_data = 12'b111011101110;
20'b00011101010111000100: color_data = 12'b111011101110;
20'b00011101010111000101: color_data = 12'b111011101110;
20'b00011101010111000110: color_data = 12'b111011101110;
20'b00011101010111000111: color_data = 12'b111011101110;
20'b00011101010111001000: color_data = 12'b111011101110;
20'b00011101010111001010: color_data = 12'b111011101110;
20'b00011101010111001011: color_data = 12'b111011101110;
20'b00011101010111001100: color_data = 12'b111011101110;
20'b00011101010111001101: color_data = 12'b111011101110;
20'b00011101010111001110: color_data = 12'b111011101110;
20'b00011101010111001111: color_data = 12'b111011101110;
20'b00011101010111010000: color_data = 12'b111011101110;
20'b00011101010111010001: color_data = 12'b111011101110;
20'b00011101010111010010: color_data = 12'b111011101110;
20'b00011101010111010011: color_data = 12'b111011101110;
20'b00011101010111010101: color_data = 12'b111011101110;
20'b00011101010111010110: color_data = 12'b111011101110;
20'b00011101010111010111: color_data = 12'b111011101110;
20'b00011101010111011000: color_data = 12'b111011101110;
20'b00011101010111011001: color_data = 12'b111011101110;
20'b00011101010111011010: color_data = 12'b111011101110;
20'b00011101010111011011: color_data = 12'b111011101110;
20'b00011101010111011100: color_data = 12'b111011101110;
20'b00011101010111011101: color_data = 12'b111011101110;
20'b00011101010111011110: color_data = 12'b111011101110;
20'b00011101010111100000: color_data = 12'b111011101110;
20'b00011101010111100001: color_data = 12'b111011101110;
20'b00011101010111100010: color_data = 12'b111011101110;
20'b00011101010111100011: color_data = 12'b111011101110;
20'b00011101010111100100: color_data = 12'b111011101110;
20'b00011101010111100101: color_data = 12'b111011101110;
20'b00011101010111100110: color_data = 12'b111011101110;
20'b00011101010111100111: color_data = 12'b111011101110;
20'b00011101010111101000: color_data = 12'b111011101110;
20'b00011101010111101001: color_data = 12'b111011101110;
20'b00011101100010101100: color_data = 12'b111011101110;
20'b00011101100010101101: color_data = 12'b111011101110;
20'b00011101100010101110: color_data = 12'b111011101110;
20'b00011101100010101111: color_data = 12'b111011101110;
20'b00011101100010110000: color_data = 12'b111011101110;
20'b00011101100010110001: color_data = 12'b111011101110;
20'b00011101100010110010: color_data = 12'b111011101110;
20'b00011101100010110011: color_data = 12'b111011101110;
20'b00011101100010110100: color_data = 12'b111011101110;
20'b00011101100010110101: color_data = 12'b111011101110;
20'b00011101100010110111: color_data = 12'b111011101110;
20'b00011101100010111000: color_data = 12'b111011101110;
20'b00011101100010111001: color_data = 12'b111011101110;
20'b00011101100010111010: color_data = 12'b111011101110;
20'b00011101100010111011: color_data = 12'b111011101110;
20'b00011101100010111100: color_data = 12'b111011101110;
20'b00011101100010111101: color_data = 12'b111011101110;
20'b00011101100010111110: color_data = 12'b111011101110;
20'b00011101100010111111: color_data = 12'b111011101110;
20'b00011101100011000000: color_data = 12'b111011101110;
20'b00011101100011000010: color_data = 12'b111011101110;
20'b00011101100011000011: color_data = 12'b111011101110;
20'b00011101100011000100: color_data = 12'b111011101110;
20'b00011101100011000101: color_data = 12'b111011101110;
20'b00011101100011000110: color_data = 12'b111011101110;
20'b00011101100011000111: color_data = 12'b111011101110;
20'b00011101100011001000: color_data = 12'b111011101110;
20'b00011101100011001001: color_data = 12'b111011101110;
20'b00011101100011001010: color_data = 12'b111011101110;
20'b00011101100011001011: color_data = 12'b111011101110;
20'b00011101100011001101: color_data = 12'b111011101110;
20'b00011101100011001110: color_data = 12'b111011101110;
20'b00011101100011001111: color_data = 12'b111011101110;
20'b00011101100011010000: color_data = 12'b111011101110;
20'b00011101100011010001: color_data = 12'b111011101110;
20'b00011101100011010010: color_data = 12'b111011101110;
20'b00011101100011010011: color_data = 12'b111011101110;
20'b00011101100011010100: color_data = 12'b111011101110;
20'b00011101100011010101: color_data = 12'b111011101110;
20'b00011101100011010110: color_data = 12'b111011101110;
20'b00011101100100000100: color_data = 12'b111011101110;
20'b00011101100100000101: color_data = 12'b111011101110;
20'b00011101100100000110: color_data = 12'b111011101110;
20'b00011101100100000111: color_data = 12'b111011101110;
20'b00011101100100001000: color_data = 12'b111011101110;
20'b00011101100100001001: color_data = 12'b111011101110;
20'b00011101100100001010: color_data = 12'b111011101110;
20'b00011101100100001011: color_data = 12'b111011101110;
20'b00011101100100001100: color_data = 12'b111011101110;
20'b00011101100100001101: color_data = 12'b111011101110;
20'b00011101100101010001: color_data = 12'b111100000000;
20'b00011101100101010010: color_data = 12'b111100000000;
20'b00011101100101010011: color_data = 12'b111100000000;
20'b00011101100101010100: color_data = 12'b111100000000;
20'b00011101100101010101: color_data = 12'b111100000000;
20'b00011101100101010110: color_data = 12'b111100000000;
20'b00011101100101010111: color_data = 12'b111100000000;
20'b00011101100101011000: color_data = 12'b111100000000;
20'b00011101100101011001: color_data = 12'b111100000000;
20'b00011101100101011010: color_data = 12'b111100000000;
20'b00011101100101011100: color_data = 12'b111100000000;
20'b00011101100101011101: color_data = 12'b111100000000;
20'b00011101100101011110: color_data = 12'b111100000000;
20'b00011101100101011111: color_data = 12'b111100000000;
20'b00011101100101100000: color_data = 12'b111100000000;
20'b00011101100101100001: color_data = 12'b111100000000;
20'b00011101100101100010: color_data = 12'b111100000000;
20'b00011101100101100011: color_data = 12'b111100000000;
20'b00011101100101100100: color_data = 12'b111100000000;
20'b00011101100101100101: color_data = 12'b111100000000;
20'b00011101100101111101: color_data = 12'b111011101110;
20'b00011101100101111110: color_data = 12'b111011101110;
20'b00011101100101111111: color_data = 12'b111011101110;
20'b00011101100110000000: color_data = 12'b111011101110;
20'b00011101100110000001: color_data = 12'b111011101110;
20'b00011101100110000010: color_data = 12'b111011101110;
20'b00011101100110000011: color_data = 12'b111011101110;
20'b00011101100110000100: color_data = 12'b111011101110;
20'b00011101100110000101: color_data = 12'b111011101110;
20'b00011101100110000110: color_data = 12'b111011101110;
20'b00011101100110001000: color_data = 12'b111011101110;
20'b00011101100110001001: color_data = 12'b111011101110;
20'b00011101100110001010: color_data = 12'b111011101110;
20'b00011101100110001011: color_data = 12'b111011101110;
20'b00011101100110001100: color_data = 12'b111011101110;
20'b00011101100110001101: color_data = 12'b111011101110;
20'b00011101100110001110: color_data = 12'b111011101110;
20'b00011101100110001111: color_data = 12'b111011101110;
20'b00011101100110010000: color_data = 12'b111011101110;
20'b00011101100110010001: color_data = 12'b111011101110;
20'b00011101100110110100: color_data = 12'b111011101110;
20'b00011101100110110101: color_data = 12'b111011101110;
20'b00011101100110110110: color_data = 12'b111011101110;
20'b00011101100110110111: color_data = 12'b111011101110;
20'b00011101100110111000: color_data = 12'b111011101110;
20'b00011101100110111001: color_data = 12'b111011101110;
20'b00011101100110111010: color_data = 12'b111011101110;
20'b00011101100110111011: color_data = 12'b111011101110;
20'b00011101100110111100: color_data = 12'b111011101110;
20'b00011101100110111101: color_data = 12'b111011101110;
20'b00011101100110111111: color_data = 12'b111011101110;
20'b00011101100111000000: color_data = 12'b111011101110;
20'b00011101100111000001: color_data = 12'b111011101110;
20'b00011101100111000010: color_data = 12'b111011101110;
20'b00011101100111000011: color_data = 12'b111011101110;
20'b00011101100111000100: color_data = 12'b111011101110;
20'b00011101100111000101: color_data = 12'b111011101110;
20'b00011101100111000110: color_data = 12'b111011101110;
20'b00011101100111000111: color_data = 12'b111011101110;
20'b00011101100111001000: color_data = 12'b111011101110;
20'b00011101100111001010: color_data = 12'b111011101110;
20'b00011101100111001011: color_data = 12'b111011101110;
20'b00011101100111001100: color_data = 12'b111011101110;
20'b00011101100111001101: color_data = 12'b111011101110;
20'b00011101100111001110: color_data = 12'b111011101110;
20'b00011101100111001111: color_data = 12'b111011101110;
20'b00011101100111010000: color_data = 12'b111011101110;
20'b00011101100111010001: color_data = 12'b111011101110;
20'b00011101100111010010: color_data = 12'b111011101110;
20'b00011101100111010011: color_data = 12'b111011101110;
20'b00011101100111010101: color_data = 12'b111011101110;
20'b00011101100111010110: color_data = 12'b111011101110;
20'b00011101100111010111: color_data = 12'b111011101110;
20'b00011101100111011000: color_data = 12'b111011101110;
20'b00011101100111011001: color_data = 12'b111011101110;
20'b00011101100111011010: color_data = 12'b111011101110;
20'b00011101100111011011: color_data = 12'b111011101110;
20'b00011101100111011100: color_data = 12'b111011101110;
20'b00011101100111011101: color_data = 12'b111011101110;
20'b00011101100111011110: color_data = 12'b111011101110;
20'b00011101100111100000: color_data = 12'b111011101110;
20'b00011101100111100001: color_data = 12'b111011101110;
20'b00011101100111100010: color_data = 12'b111011101110;
20'b00011101100111100011: color_data = 12'b111011101110;
20'b00011101100111100100: color_data = 12'b111011101110;
20'b00011101100111100101: color_data = 12'b111011101110;
20'b00011101100111100110: color_data = 12'b111011101110;
20'b00011101100111100111: color_data = 12'b111011101110;
20'b00011101100111101000: color_data = 12'b111011101110;
20'b00011101100111101001: color_data = 12'b111011101110;
20'b00011101110010101100: color_data = 12'b111011101110;
20'b00011101110010101101: color_data = 12'b111011101110;
20'b00011101110010101110: color_data = 12'b111011101110;
20'b00011101110010101111: color_data = 12'b111011101110;
20'b00011101110010110000: color_data = 12'b111011101110;
20'b00011101110010110001: color_data = 12'b111011101110;
20'b00011101110010110010: color_data = 12'b111011101110;
20'b00011101110010110011: color_data = 12'b111011101110;
20'b00011101110010110100: color_data = 12'b111011101110;
20'b00011101110010110101: color_data = 12'b111011101110;
20'b00011101110010110111: color_data = 12'b111011101110;
20'b00011101110010111000: color_data = 12'b111011101110;
20'b00011101110010111001: color_data = 12'b111011101110;
20'b00011101110010111010: color_data = 12'b111011101110;
20'b00011101110010111011: color_data = 12'b111011101110;
20'b00011101110010111100: color_data = 12'b111011101110;
20'b00011101110010111101: color_data = 12'b111011101110;
20'b00011101110010111110: color_data = 12'b111011101110;
20'b00011101110010111111: color_data = 12'b111011101110;
20'b00011101110011000000: color_data = 12'b111011101110;
20'b00011101110011000010: color_data = 12'b111011101110;
20'b00011101110011000011: color_data = 12'b111011101110;
20'b00011101110011000100: color_data = 12'b111011101110;
20'b00011101110011000101: color_data = 12'b111011101110;
20'b00011101110011000110: color_data = 12'b111011101110;
20'b00011101110011000111: color_data = 12'b111011101110;
20'b00011101110011001000: color_data = 12'b111011101110;
20'b00011101110011001001: color_data = 12'b111011101110;
20'b00011101110011001010: color_data = 12'b111011101110;
20'b00011101110011001011: color_data = 12'b111011101110;
20'b00011101110011001101: color_data = 12'b111011101110;
20'b00011101110011001110: color_data = 12'b111011101110;
20'b00011101110011001111: color_data = 12'b111011101110;
20'b00011101110011010000: color_data = 12'b111011101110;
20'b00011101110011010001: color_data = 12'b111011101110;
20'b00011101110011010010: color_data = 12'b111011101110;
20'b00011101110011010011: color_data = 12'b111011101110;
20'b00011101110011010100: color_data = 12'b111011101110;
20'b00011101110011010101: color_data = 12'b111011101110;
20'b00011101110011010110: color_data = 12'b111011101110;
20'b00011101110100000100: color_data = 12'b111011101110;
20'b00011101110100000101: color_data = 12'b111011101110;
20'b00011101110100000110: color_data = 12'b111011101110;
20'b00011101110100000111: color_data = 12'b111011101110;
20'b00011101110100001000: color_data = 12'b111011101110;
20'b00011101110100001001: color_data = 12'b111011101110;
20'b00011101110100001010: color_data = 12'b111011101110;
20'b00011101110100001011: color_data = 12'b111011101110;
20'b00011101110100001100: color_data = 12'b111011101110;
20'b00011101110100001101: color_data = 12'b111011101110;
20'b00011101110101010001: color_data = 12'b111100000000;
20'b00011101110101010010: color_data = 12'b111100000000;
20'b00011101110101010011: color_data = 12'b111100000000;
20'b00011101110101010100: color_data = 12'b111100000000;
20'b00011101110101010101: color_data = 12'b111100000000;
20'b00011101110101010110: color_data = 12'b111100000000;
20'b00011101110101010111: color_data = 12'b111100000000;
20'b00011101110101011000: color_data = 12'b111100000000;
20'b00011101110101011001: color_data = 12'b111100000000;
20'b00011101110101011010: color_data = 12'b111100000000;
20'b00011101110101011100: color_data = 12'b111100000000;
20'b00011101110101011101: color_data = 12'b111100000000;
20'b00011101110101011110: color_data = 12'b111100000000;
20'b00011101110101011111: color_data = 12'b111100000000;
20'b00011101110101100000: color_data = 12'b111100000000;
20'b00011101110101100001: color_data = 12'b111100000000;
20'b00011101110101100010: color_data = 12'b111100000000;
20'b00011101110101100011: color_data = 12'b111100000000;
20'b00011101110101100100: color_data = 12'b111100000000;
20'b00011101110101100101: color_data = 12'b111100000000;
20'b00011101110101111101: color_data = 12'b111011101110;
20'b00011101110101111110: color_data = 12'b111011101110;
20'b00011101110101111111: color_data = 12'b111011101110;
20'b00011101110110000000: color_data = 12'b111011101110;
20'b00011101110110000001: color_data = 12'b111011101110;
20'b00011101110110000010: color_data = 12'b111011101110;
20'b00011101110110000011: color_data = 12'b111011101110;
20'b00011101110110000100: color_data = 12'b111011101110;
20'b00011101110110000101: color_data = 12'b111011101110;
20'b00011101110110000110: color_data = 12'b111011101110;
20'b00011101110110001000: color_data = 12'b111011101110;
20'b00011101110110001001: color_data = 12'b111011101110;
20'b00011101110110001010: color_data = 12'b111011101110;
20'b00011101110110001011: color_data = 12'b111011101110;
20'b00011101110110001100: color_data = 12'b111011101110;
20'b00011101110110001101: color_data = 12'b111011101110;
20'b00011101110110001110: color_data = 12'b111011101110;
20'b00011101110110001111: color_data = 12'b111011101110;
20'b00011101110110010000: color_data = 12'b111011101110;
20'b00011101110110010001: color_data = 12'b111011101110;
20'b00011101110110110100: color_data = 12'b111011101110;
20'b00011101110110110101: color_data = 12'b111011101110;
20'b00011101110110110110: color_data = 12'b111011101110;
20'b00011101110110110111: color_data = 12'b111011101110;
20'b00011101110110111000: color_data = 12'b111011101110;
20'b00011101110110111001: color_data = 12'b111011101110;
20'b00011101110110111010: color_data = 12'b111011101110;
20'b00011101110110111011: color_data = 12'b111011101110;
20'b00011101110110111100: color_data = 12'b111011101110;
20'b00011101110110111101: color_data = 12'b111011101110;
20'b00011101110110111111: color_data = 12'b111011101110;
20'b00011101110111000000: color_data = 12'b111011101110;
20'b00011101110111000001: color_data = 12'b111011101110;
20'b00011101110111000010: color_data = 12'b111011101110;
20'b00011101110111000011: color_data = 12'b111011101110;
20'b00011101110111000100: color_data = 12'b111011101110;
20'b00011101110111000101: color_data = 12'b111011101110;
20'b00011101110111000110: color_data = 12'b111011101110;
20'b00011101110111000111: color_data = 12'b111011101110;
20'b00011101110111001000: color_data = 12'b111011101110;
20'b00011101110111001010: color_data = 12'b111011101110;
20'b00011101110111001011: color_data = 12'b111011101110;
20'b00011101110111001100: color_data = 12'b111011101110;
20'b00011101110111001101: color_data = 12'b111011101110;
20'b00011101110111001110: color_data = 12'b111011101110;
20'b00011101110111001111: color_data = 12'b111011101110;
20'b00011101110111010000: color_data = 12'b111011101110;
20'b00011101110111010001: color_data = 12'b111011101110;
20'b00011101110111010010: color_data = 12'b111011101110;
20'b00011101110111010011: color_data = 12'b111011101110;
20'b00011101110111010101: color_data = 12'b111011101110;
20'b00011101110111010110: color_data = 12'b111011101110;
20'b00011101110111010111: color_data = 12'b111011101110;
20'b00011101110111011000: color_data = 12'b111011101110;
20'b00011101110111011001: color_data = 12'b111011101110;
20'b00011101110111011010: color_data = 12'b111011101110;
20'b00011101110111011011: color_data = 12'b111011101110;
20'b00011101110111011100: color_data = 12'b111011101110;
20'b00011101110111011101: color_data = 12'b111011101110;
20'b00011101110111011110: color_data = 12'b111011101110;
20'b00011101110111100000: color_data = 12'b111011101110;
20'b00011101110111100001: color_data = 12'b111011101110;
20'b00011101110111100010: color_data = 12'b111011101110;
20'b00011101110111100011: color_data = 12'b111011101110;
20'b00011101110111100100: color_data = 12'b111011101110;
20'b00011101110111100101: color_data = 12'b111011101110;
20'b00011101110111100110: color_data = 12'b111011101110;
20'b00011101110111100111: color_data = 12'b111011101110;
20'b00011101110111101000: color_data = 12'b111011101110;
20'b00011101110111101001: color_data = 12'b111011101110;
20'b00011110000010101100: color_data = 12'b111011101110;
20'b00011110000010101101: color_data = 12'b111011101110;
20'b00011110000010101110: color_data = 12'b111011101110;
20'b00011110000010101111: color_data = 12'b111011101110;
20'b00011110000010110000: color_data = 12'b111011101110;
20'b00011110000010110001: color_data = 12'b111011101110;
20'b00011110000010110010: color_data = 12'b111011101110;
20'b00011110000010110011: color_data = 12'b111011101110;
20'b00011110000010110100: color_data = 12'b111011101110;
20'b00011110000010110101: color_data = 12'b111011101110;
20'b00011110000010110111: color_data = 12'b111011101110;
20'b00011110000010111000: color_data = 12'b111011101110;
20'b00011110000010111001: color_data = 12'b111011101110;
20'b00011110000010111010: color_data = 12'b111011101110;
20'b00011110000010111011: color_data = 12'b111011101110;
20'b00011110000010111100: color_data = 12'b111011101110;
20'b00011110000010111101: color_data = 12'b111011101110;
20'b00011110000010111110: color_data = 12'b111011101110;
20'b00011110000010111111: color_data = 12'b111011101110;
20'b00011110000011000000: color_data = 12'b111011101110;
20'b00011110000011000010: color_data = 12'b111011101110;
20'b00011110000011000011: color_data = 12'b111011101110;
20'b00011110000011000100: color_data = 12'b111011101110;
20'b00011110000011000101: color_data = 12'b111011101110;
20'b00011110000011000110: color_data = 12'b111011101110;
20'b00011110000011000111: color_data = 12'b111011101110;
20'b00011110000011001000: color_data = 12'b111011101110;
20'b00011110000011001001: color_data = 12'b111011101110;
20'b00011110000011001010: color_data = 12'b111011101110;
20'b00011110000011001011: color_data = 12'b111011101110;
20'b00011110000011001101: color_data = 12'b111011101110;
20'b00011110000011001110: color_data = 12'b111011101110;
20'b00011110000011001111: color_data = 12'b111011101110;
20'b00011110000011010000: color_data = 12'b111011101110;
20'b00011110000011010001: color_data = 12'b111011101110;
20'b00011110000011010010: color_data = 12'b111011101110;
20'b00011110000011010011: color_data = 12'b111011101110;
20'b00011110000011010100: color_data = 12'b111011101110;
20'b00011110000011010101: color_data = 12'b111011101110;
20'b00011110000011010110: color_data = 12'b111011101110;
20'b00011110000100000100: color_data = 12'b111011101110;
20'b00011110000100000101: color_data = 12'b111011101110;
20'b00011110000100000110: color_data = 12'b111011101110;
20'b00011110000100000111: color_data = 12'b111011101110;
20'b00011110000100001000: color_data = 12'b111011101110;
20'b00011110000100001001: color_data = 12'b111011101110;
20'b00011110000100001010: color_data = 12'b111011101110;
20'b00011110000100001011: color_data = 12'b111011101110;
20'b00011110000100001100: color_data = 12'b111011101110;
20'b00011110000100001101: color_data = 12'b111011101110;
20'b00011110000101010001: color_data = 12'b111100000000;
20'b00011110000101010010: color_data = 12'b111100000000;
20'b00011110000101010011: color_data = 12'b111100000000;
20'b00011110000101010100: color_data = 12'b111100000000;
20'b00011110000101010101: color_data = 12'b111100000000;
20'b00011110000101010110: color_data = 12'b111100000000;
20'b00011110000101010111: color_data = 12'b111100000000;
20'b00011110000101011000: color_data = 12'b111100000000;
20'b00011110000101011001: color_data = 12'b111100000000;
20'b00011110000101011010: color_data = 12'b111100000000;
20'b00011110000101011100: color_data = 12'b111100000000;
20'b00011110000101011101: color_data = 12'b111100000000;
20'b00011110000101011110: color_data = 12'b111100000000;
20'b00011110000101011111: color_data = 12'b111100000000;
20'b00011110000101100000: color_data = 12'b111100000000;
20'b00011110000101100001: color_data = 12'b111100000000;
20'b00011110000101100010: color_data = 12'b111100000000;
20'b00011110000101100011: color_data = 12'b111100000000;
20'b00011110000101100100: color_data = 12'b111100000000;
20'b00011110000101100101: color_data = 12'b111100000000;
20'b00011110000101111101: color_data = 12'b111011101110;
20'b00011110000101111110: color_data = 12'b111011101110;
20'b00011110000101111111: color_data = 12'b111011101110;
20'b00011110000110000000: color_data = 12'b111011101110;
20'b00011110000110000001: color_data = 12'b111011101110;
20'b00011110000110000010: color_data = 12'b111011101110;
20'b00011110000110000011: color_data = 12'b111011101110;
20'b00011110000110000100: color_data = 12'b111011101110;
20'b00011110000110000101: color_data = 12'b111011101110;
20'b00011110000110000110: color_data = 12'b111011101110;
20'b00011110000110001000: color_data = 12'b111011101110;
20'b00011110000110001001: color_data = 12'b111011101110;
20'b00011110000110001010: color_data = 12'b111011101110;
20'b00011110000110001011: color_data = 12'b111011101110;
20'b00011110000110001100: color_data = 12'b111011101110;
20'b00011110000110001101: color_data = 12'b111011101110;
20'b00011110000110001110: color_data = 12'b111011101110;
20'b00011110000110001111: color_data = 12'b111011101110;
20'b00011110000110010000: color_data = 12'b111011101110;
20'b00011110000110010001: color_data = 12'b111011101110;
20'b00011110000110110100: color_data = 12'b111011101110;
20'b00011110000110110101: color_data = 12'b111011101110;
20'b00011110000110110110: color_data = 12'b111011101110;
20'b00011110000110110111: color_data = 12'b111011101110;
20'b00011110000110111000: color_data = 12'b111011101110;
20'b00011110000110111001: color_data = 12'b111011101110;
20'b00011110000110111010: color_data = 12'b111011101110;
20'b00011110000110111011: color_data = 12'b111011101110;
20'b00011110000110111100: color_data = 12'b111011101110;
20'b00011110000110111101: color_data = 12'b111011101110;
20'b00011110000110111111: color_data = 12'b111011101110;
20'b00011110000111000000: color_data = 12'b111011101110;
20'b00011110000111000001: color_data = 12'b111011101110;
20'b00011110000111000010: color_data = 12'b111011101110;
20'b00011110000111000011: color_data = 12'b111011101110;
20'b00011110000111000100: color_data = 12'b111011101110;
20'b00011110000111000101: color_data = 12'b111011101110;
20'b00011110000111000110: color_data = 12'b111011101110;
20'b00011110000111000111: color_data = 12'b111011101110;
20'b00011110000111001000: color_data = 12'b111011101110;
20'b00011110000111001010: color_data = 12'b111011101110;
20'b00011110000111001011: color_data = 12'b111011101110;
20'b00011110000111001100: color_data = 12'b111011101110;
20'b00011110000111001101: color_data = 12'b111011101110;
20'b00011110000111001110: color_data = 12'b111011101110;
20'b00011110000111001111: color_data = 12'b111011101110;
20'b00011110000111010000: color_data = 12'b111011101110;
20'b00011110000111010001: color_data = 12'b111011101110;
20'b00011110000111010010: color_data = 12'b111011101110;
20'b00011110000111010011: color_data = 12'b111011101110;
20'b00011110000111010101: color_data = 12'b111011101110;
20'b00011110000111010110: color_data = 12'b111011101110;
20'b00011110000111010111: color_data = 12'b111011101110;
20'b00011110000111011000: color_data = 12'b111011101110;
20'b00011110000111011001: color_data = 12'b111011101110;
20'b00011110000111011010: color_data = 12'b111011101110;
20'b00011110000111011011: color_data = 12'b111011101110;
20'b00011110000111011100: color_data = 12'b111011101110;
20'b00011110000111011101: color_data = 12'b111011101110;
20'b00011110000111011110: color_data = 12'b111011101110;
20'b00011110000111100000: color_data = 12'b111011101110;
20'b00011110000111100001: color_data = 12'b111011101110;
20'b00011110000111100010: color_data = 12'b111011101110;
20'b00011110000111100011: color_data = 12'b111011101110;
20'b00011110000111100100: color_data = 12'b111011101110;
20'b00011110000111100101: color_data = 12'b111011101110;
20'b00011110000111100110: color_data = 12'b111011101110;
20'b00011110000111100111: color_data = 12'b111011101110;
20'b00011110000111101000: color_data = 12'b111011101110;
20'b00011110000111101001: color_data = 12'b111011101110;
20'b00011110010010101100: color_data = 12'b111011101110;
20'b00011110010010101101: color_data = 12'b111011101110;
20'b00011110010010101110: color_data = 12'b111011101110;
20'b00011110010010101111: color_data = 12'b111011101110;
20'b00011110010010110000: color_data = 12'b111011101110;
20'b00011110010010110001: color_data = 12'b111011101110;
20'b00011110010010110010: color_data = 12'b111011101110;
20'b00011110010010110011: color_data = 12'b111011101110;
20'b00011110010010110100: color_data = 12'b111011101110;
20'b00011110010010110101: color_data = 12'b111011101110;
20'b00011110010010110111: color_data = 12'b111011101110;
20'b00011110010010111000: color_data = 12'b111011101110;
20'b00011110010010111001: color_data = 12'b111011101110;
20'b00011110010010111010: color_data = 12'b111011101110;
20'b00011110010010111011: color_data = 12'b111011101110;
20'b00011110010010111100: color_data = 12'b111011101110;
20'b00011110010010111101: color_data = 12'b111011101110;
20'b00011110010010111110: color_data = 12'b111011101110;
20'b00011110010010111111: color_data = 12'b111011101110;
20'b00011110010011000000: color_data = 12'b111011101110;
20'b00011110010011000010: color_data = 12'b111011101110;
20'b00011110010011000011: color_data = 12'b111011101110;
20'b00011110010011000100: color_data = 12'b111011101110;
20'b00011110010011000101: color_data = 12'b111011101110;
20'b00011110010011000110: color_data = 12'b111011101110;
20'b00011110010011000111: color_data = 12'b111011101110;
20'b00011110010011001000: color_data = 12'b111011101110;
20'b00011110010011001001: color_data = 12'b111011101110;
20'b00011110010011001010: color_data = 12'b111011101110;
20'b00011110010011001011: color_data = 12'b111011101110;
20'b00011110010011001101: color_data = 12'b111011101110;
20'b00011110010011001110: color_data = 12'b111011101110;
20'b00011110010011001111: color_data = 12'b111011101110;
20'b00011110010011010000: color_data = 12'b111011101110;
20'b00011110010011010001: color_data = 12'b111011101110;
20'b00011110010011010010: color_data = 12'b111011101110;
20'b00011110010011010011: color_data = 12'b111011101110;
20'b00011110010011010100: color_data = 12'b111011101110;
20'b00011110010011010101: color_data = 12'b111011101110;
20'b00011110010011010110: color_data = 12'b111011101110;
20'b00011110010100000100: color_data = 12'b111011101110;
20'b00011110010100000101: color_data = 12'b111011101110;
20'b00011110010100000110: color_data = 12'b111011101110;
20'b00011110010100000111: color_data = 12'b111011101110;
20'b00011110010100001000: color_data = 12'b111011101110;
20'b00011110010100001001: color_data = 12'b111011101110;
20'b00011110010100001010: color_data = 12'b111011101110;
20'b00011110010100001011: color_data = 12'b111011101110;
20'b00011110010100001100: color_data = 12'b111011101110;
20'b00011110010100001101: color_data = 12'b111011101110;
20'b00011110010101010001: color_data = 12'b111100000000;
20'b00011110010101010010: color_data = 12'b111100000000;
20'b00011110010101010011: color_data = 12'b111100000000;
20'b00011110010101010100: color_data = 12'b111100000000;
20'b00011110010101010101: color_data = 12'b111100000000;
20'b00011110010101010110: color_data = 12'b111100000000;
20'b00011110010101010111: color_data = 12'b111100000000;
20'b00011110010101011000: color_data = 12'b111100000000;
20'b00011110010101011001: color_data = 12'b111100000000;
20'b00011110010101011010: color_data = 12'b111100000000;
20'b00011110010101011100: color_data = 12'b111100000000;
20'b00011110010101011101: color_data = 12'b111100000000;
20'b00011110010101011110: color_data = 12'b111100000000;
20'b00011110010101011111: color_data = 12'b111100000000;
20'b00011110010101100000: color_data = 12'b111100000000;
20'b00011110010101100001: color_data = 12'b111100000000;
20'b00011110010101100010: color_data = 12'b111100000000;
20'b00011110010101100011: color_data = 12'b111100000000;
20'b00011110010101100100: color_data = 12'b111100000000;
20'b00011110010101100101: color_data = 12'b111100000000;
20'b00011110010101111101: color_data = 12'b111011101110;
20'b00011110010101111110: color_data = 12'b111011101110;
20'b00011110010101111111: color_data = 12'b111011101110;
20'b00011110010110000000: color_data = 12'b111011101110;
20'b00011110010110000001: color_data = 12'b111011101110;
20'b00011110010110000010: color_data = 12'b111011101110;
20'b00011110010110000011: color_data = 12'b111011101110;
20'b00011110010110000100: color_data = 12'b111011101110;
20'b00011110010110000101: color_data = 12'b111011101110;
20'b00011110010110000110: color_data = 12'b111011101110;
20'b00011110010110001000: color_data = 12'b111011101110;
20'b00011110010110001001: color_data = 12'b111011101110;
20'b00011110010110001010: color_data = 12'b111011101110;
20'b00011110010110001011: color_data = 12'b111011101110;
20'b00011110010110001100: color_data = 12'b111011101110;
20'b00011110010110001101: color_data = 12'b111011101110;
20'b00011110010110001110: color_data = 12'b111011101110;
20'b00011110010110001111: color_data = 12'b111011101110;
20'b00011110010110010000: color_data = 12'b111011101110;
20'b00011110010110010001: color_data = 12'b111011101110;
20'b00011110010110110100: color_data = 12'b111011101110;
20'b00011110010110110101: color_data = 12'b111011101110;
20'b00011110010110110110: color_data = 12'b111011101110;
20'b00011110010110110111: color_data = 12'b111011101110;
20'b00011110010110111000: color_data = 12'b111011101110;
20'b00011110010110111001: color_data = 12'b111011101110;
20'b00011110010110111010: color_data = 12'b111011101110;
20'b00011110010110111011: color_data = 12'b111011101110;
20'b00011110010110111100: color_data = 12'b111011101110;
20'b00011110010110111101: color_data = 12'b111011101110;
20'b00011110010110111111: color_data = 12'b111011101110;
20'b00011110010111000000: color_data = 12'b111011101110;
20'b00011110010111000001: color_data = 12'b111011101110;
20'b00011110010111000010: color_data = 12'b111011101110;
20'b00011110010111000011: color_data = 12'b111011101110;
20'b00011110010111000100: color_data = 12'b111011101110;
20'b00011110010111000101: color_data = 12'b111011101110;
20'b00011110010111000110: color_data = 12'b111011101110;
20'b00011110010111000111: color_data = 12'b111011101110;
20'b00011110010111001000: color_data = 12'b111011101110;
20'b00011110010111001010: color_data = 12'b111011101110;
20'b00011110010111001011: color_data = 12'b111011101110;
20'b00011110010111001100: color_data = 12'b111011101110;
20'b00011110010111001101: color_data = 12'b111011101110;
20'b00011110010111001110: color_data = 12'b111011101110;
20'b00011110010111001111: color_data = 12'b111011101110;
20'b00011110010111010000: color_data = 12'b111011101110;
20'b00011110010111010001: color_data = 12'b111011101110;
20'b00011110010111010010: color_data = 12'b111011101110;
20'b00011110010111010011: color_data = 12'b111011101110;
20'b00011110010111010101: color_data = 12'b111011101110;
20'b00011110010111010110: color_data = 12'b111011101110;
20'b00011110010111010111: color_data = 12'b111011101110;
20'b00011110010111011000: color_data = 12'b111011101110;
20'b00011110010111011001: color_data = 12'b111011101110;
20'b00011110010111011010: color_data = 12'b111011101110;
20'b00011110010111011011: color_data = 12'b111011101110;
20'b00011110010111011100: color_data = 12'b111011101110;
20'b00011110010111011101: color_data = 12'b111011101110;
20'b00011110010111011110: color_data = 12'b111011101110;
20'b00011110010111100000: color_data = 12'b111011101110;
20'b00011110010111100001: color_data = 12'b111011101110;
20'b00011110010111100010: color_data = 12'b111011101110;
20'b00011110010111100011: color_data = 12'b111011101110;
20'b00011110010111100100: color_data = 12'b111011101110;
20'b00011110010111100101: color_data = 12'b111011101110;
20'b00011110010111100110: color_data = 12'b111011101110;
20'b00011110010111100111: color_data = 12'b111011101110;
20'b00011110010111101000: color_data = 12'b111011101110;
20'b00011110010111101001: color_data = 12'b111011101110;
20'b00011110100010101100: color_data = 12'b111011101110;
20'b00011110100010101101: color_data = 12'b111011101110;
20'b00011110100010101110: color_data = 12'b111011101110;
20'b00011110100010101111: color_data = 12'b111011101110;
20'b00011110100010110000: color_data = 12'b111011101110;
20'b00011110100010110001: color_data = 12'b111011101110;
20'b00011110100010110010: color_data = 12'b111011101110;
20'b00011110100010110011: color_data = 12'b111011101110;
20'b00011110100010110100: color_data = 12'b111011101110;
20'b00011110100010110101: color_data = 12'b111011101110;
20'b00011110100010110111: color_data = 12'b111011101110;
20'b00011110100010111000: color_data = 12'b111011101110;
20'b00011110100010111001: color_data = 12'b111011101110;
20'b00011110100010111010: color_data = 12'b111011101110;
20'b00011110100010111011: color_data = 12'b111011101110;
20'b00011110100010111100: color_data = 12'b111011101110;
20'b00011110100010111101: color_data = 12'b111011101110;
20'b00011110100010111110: color_data = 12'b111011101110;
20'b00011110100010111111: color_data = 12'b111011101110;
20'b00011110100011000000: color_data = 12'b111011101110;
20'b00011110100011000010: color_data = 12'b111011101110;
20'b00011110100011000011: color_data = 12'b111011101110;
20'b00011110100011000100: color_data = 12'b111011101110;
20'b00011110100011000101: color_data = 12'b111011101110;
20'b00011110100011000110: color_data = 12'b111011101110;
20'b00011110100011000111: color_data = 12'b111011101110;
20'b00011110100011001000: color_data = 12'b111011101110;
20'b00011110100011001001: color_data = 12'b111011101110;
20'b00011110100011001010: color_data = 12'b111011101110;
20'b00011110100011001011: color_data = 12'b111011101110;
20'b00011110100011001101: color_data = 12'b111011101110;
20'b00011110100011001110: color_data = 12'b111011101110;
20'b00011110100011001111: color_data = 12'b111011101110;
20'b00011110100011010000: color_data = 12'b111011101110;
20'b00011110100011010001: color_data = 12'b111011101110;
20'b00011110100011010010: color_data = 12'b111011101110;
20'b00011110100011010011: color_data = 12'b111011101110;
20'b00011110100011010100: color_data = 12'b111011101110;
20'b00011110100011010101: color_data = 12'b111011101110;
20'b00011110100011010110: color_data = 12'b111011101110;
20'b00011110100100000100: color_data = 12'b111011101110;
20'b00011110100100000101: color_data = 12'b111011101110;
20'b00011110100100000110: color_data = 12'b111011101110;
20'b00011110100100000111: color_data = 12'b111011101110;
20'b00011110100100001000: color_data = 12'b111011101110;
20'b00011110100100001001: color_data = 12'b111011101110;
20'b00011110100100001010: color_data = 12'b111011101110;
20'b00011110100100001011: color_data = 12'b111011101110;
20'b00011110100100001100: color_data = 12'b111011101110;
20'b00011110100100001101: color_data = 12'b111011101110;
20'b00011110100101010001: color_data = 12'b111100000000;
20'b00011110100101010010: color_data = 12'b111100000000;
20'b00011110100101010011: color_data = 12'b111100000000;
20'b00011110100101010100: color_data = 12'b111100000000;
20'b00011110100101010101: color_data = 12'b111100000000;
20'b00011110100101010110: color_data = 12'b111100000000;
20'b00011110100101010111: color_data = 12'b111100000000;
20'b00011110100101011000: color_data = 12'b111100000000;
20'b00011110100101011001: color_data = 12'b111100000000;
20'b00011110100101011010: color_data = 12'b111100000000;
20'b00011110100101011100: color_data = 12'b111100000000;
20'b00011110100101011101: color_data = 12'b111100000000;
20'b00011110100101011110: color_data = 12'b111100000000;
20'b00011110100101011111: color_data = 12'b111100000000;
20'b00011110100101100000: color_data = 12'b111100000000;
20'b00011110100101100001: color_data = 12'b111100000000;
20'b00011110100101100010: color_data = 12'b111100000000;
20'b00011110100101100011: color_data = 12'b111100000000;
20'b00011110100101100100: color_data = 12'b111100000000;
20'b00011110100101100101: color_data = 12'b111100000000;
20'b00011110100101111101: color_data = 12'b111011101110;
20'b00011110100101111110: color_data = 12'b111011101110;
20'b00011110100101111111: color_data = 12'b111011101110;
20'b00011110100110000000: color_data = 12'b111011101110;
20'b00011110100110000001: color_data = 12'b111011101110;
20'b00011110100110000010: color_data = 12'b111011101110;
20'b00011110100110000011: color_data = 12'b111011101110;
20'b00011110100110000100: color_data = 12'b111011101110;
20'b00011110100110000101: color_data = 12'b111011101110;
20'b00011110100110000110: color_data = 12'b111011101110;
20'b00011110100110001000: color_data = 12'b111011101110;
20'b00011110100110001001: color_data = 12'b111011101110;
20'b00011110100110001010: color_data = 12'b111011101110;
20'b00011110100110001011: color_data = 12'b111011101110;
20'b00011110100110001100: color_data = 12'b111011101110;
20'b00011110100110001101: color_data = 12'b111011101110;
20'b00011110100110001110: color_data = 12'b111011101110;
20'b00011110100110001111: color_data = 12'b111011101110;
20'b00011110100110010000: color_data = 12'b111011101110;
20'b00011110100110010001: color_data = 12'b111011101110;
20'b00011110100110110100: color_data = 12'b111011101110;
20'b00011110100110110101: color_data = 12'b111011101110;
20'b00011110100110110110: color_data = 12'b111011101110;
20'b00011110100110110111: color_data = 12'b111011101110;
20'b00011110100110111000: color_data = 12'b111011101110;
20'b00011110100110111001: color_data = 12'b111011101110;
20'b00011110100110111010: color_data = 12'b111011101110;
20'b00011110100110111011: color_data = 12'b111011101110;
20'b00011110100110111100: color_data = 12'b111011101110;
20'b00011110100110111101: color_data = 12'b111011101110;
20'b00011110100110111111: color_data = 12'b111011101110;
20'b00011110100111000000: color_data = 12'b111011101110;
20'b00011110100111000001: color_data = 12'b111011101110;
20'b00011110100111000010: color_data = 12'b111011101110;
20'b00011110100111000011: color_data = 12'b111011101110;
20'b00011110100111000100: color_data = 12'b111011101110;
20'b00011110100111000101: color_data = 12'b111011101110;
20'b00011110100111000110: color_data = 12'b111011101110;
20'b00011110100111000111: color_data = 12'b111011101110;
20'b00011110100111001000: color_data = 12'b111011101110;
20'b00011110100111001010: color_data = 12'b111011101110;
20'b00011110100111001011: color_data = 12'b111011101110;
20'b00011110100111001100: color_data = 12'b111011101110;
20'b00011110100111001101: color_data = 12'b111011101110;
20'b00011110100111001110: color_data = 12'b111011101110;
20'b00011110100111001111: color_data = 12'b111011101110;
20'b00011110100111010000: color_data = 12'b111011101110;
20'b00011110100111010001: color_data = 12'b111011101110;
20'b00011110100111010010: color_data = 12'b111011101110;
20'b00011110100111010011: color_data = 12'b111011101110;
20'b00011110100111010101: color_data = 12'b111011101110;
20'b00011110100111010110: color_data = 12'b111011101110;
20'b00011110100111010111: color_data = 12'b111011101110;
20'b00011110100111011000: color_data = 12'b111011101110;
20'b00011110100111011001: color_data = 12'b111011101110;
20'b00011110100111011010: color_data = 12'b111011101110;
20'b00011110100111011011: color_data = 12'b111011101110;
20'b00011110100111011100: color_data = 12'b111011101110;
20'b00011110100111011101: color_data = 12'b111011101110;
20'b00011110100111011110: color_data = 12'b111011101110;
20'b00011110100111100000: color_data = 12'b111011101110;
20'b00011110100111100001: color_data = 12'b111011101110;
20'b00011110100111100010: color_data = 12'b111011101110;
20'b00011110100111100011: color_data = 12'b111011101110;
20'b00011110100111100100: color_data = 12'b111011101110;
20'b00011110100111100101: color_data = 12'b111011101110;
20'b00011110100111100110: color_data = 12'b111011101110;
20'b00011110100111100111: color_data = 12'b111011101110;
20'b00011110100111101000: color_data = 12'b111011101110;
20'b00011110100111101001: color_data = 12'b111011101110;
20'b00011110110010101100: color_data = 12'b111011101110;
20'b00011110110010101101: color_data = 12'b111011101110;
20'b00011110110010101110: color_data = 12'b111011101110;
20'b00011110110010101111: color_data = 12'b111011101110;
20'b00011110110010110000: color_data = 12'b111011101110;
20'b00011110110010110001: color_data = 12'b111011101110;
20'b00011110110010110010: color_data = 12'b111011101110;
20'b00011110110010110011: color_data = 12'b111011101110;
20'b00011110110010110100: color_data = 12'b111011101110;
20'b00011110110010110101: color_data = 12'b111011101110;
20'b00011110110010110111: color_data = 12'b111011101110;
20'b00011110110010111000: color_data = 12'b111011101110;
20'b00011110110010111001: color_data = 12'b111011101110;
20'b00011110110010111010: color_data = 12'b111011101110;
20'b00011110110010111011: color_data = 12'b111011101110;
20'b00011110110010111100: color_data = 12'b111011101110;
20'b00011110110010111101: color_data = 12'b111011101110;
20'b00011110110010111110: color_data = 12'b111011101110;
20'b00011110110010111111: color_data = 12'b111011101110;
20'b00011110110011000000: color_data = 12'b111011101110;
20'b00011110110011000010: color_data = 12'b111011101110;
20'b00011110110011000011: color_data = 12'b111011101110;
20'b00011110110011000100: color_data = 12'b111011101110;
20'b00011110110011000101: color_data = 12'b111011101110;
20'b00011110110011000110: color_data = 12'b111011101110;
20'b00011110110011000111: color_data = 12'b111011101110;
20'b00011110110011001000: color_data = 12'b111011101110;
20'b00011110110011001001: color_data = 12'b111011101110;
20'b00011110110011001010: color_data = 12'b111011101110;
20'b00011110110011001011: color_data = 12'b111011101110;
20'b00011110110011001101: color_data = 12'b111011101110;
20'b00011110110011001110: color_data = 12'b111011101110;
20'b00011110110011001111: color_data = 12'b111011101110;
20'b00011110110011010000: color_data = 12'b111011101110;
20'b00011110110011010001: color_data = 12'b111011101110;
20'b00011110110011010010: color_data = 12'b111011101110;
20'b00011110110011010011: color_data = 12'b111011101110;
20'b00011110110011010100: color_data = 12'b111011101110;
20'b00011110110011010101: color_data = 12'b111011101110;
20'b00011110110011010110: color_data = 12'b111011101110;
20'b00011110110100000100: color_data = 12'b111011101110;
20'b00011110110100000101: color_data = 12'b111011101110;
20'b00011110110100000110: color_data = 12'b111011101110;
20'b00011110110100000111: color_data = 12'b111011101110;
20'b00011110110100001000: color_data = 12'b111011101110;
20'b00011110110100001001: color_data = 12'b111011101110;
20'b00011110110100001010: color_data = 12'b111011101110;
20'b00011110110100001011: color_data = 12'b111011101110;
20'b00011110110100001100: color_data = 12'b111011101110;
20'b00011110110100001101: color_data = 12'b111011101110;
20'b00011110110101010001: color_data = 12'b111100000000;
20'b00011110110101010010: color_data = 12'b111100000000;
20'b00011110110101010011: color_data = 12'b111100000000;
20'b00011110110101010100: color_data = 12'b111100000000;
20'b00011110110101010101: color_data = 12'b111100000000;
20'b00011110110101010110: color_data = 12'b111100000000;
20'b00011110110101010111: color_data = 12'b111100000000;
20'b00011110110101011000: color_data = 12'b111100000000;
20'b00011110110101011001: color_data = 12'b111100000000;
20'b00011110110101011010: color_data = 12'b111100000000;
20'b00011110110101011100: color_data = 12'b111100000000;
20'b00011110110101011101: color_data = 12'b111100000000;
20'b00011110110101011110: color_data = 12'b111100000000;
20'b00011110110101011111: color_data = 12'b111100000000;
20'b00011110110101100000: color_data = 12'b111100000000;
20'b00011110110101100001: color_data = 12'b111100000000;
20'b00011110110101100010: color_data = 12'b111100000000;
20'b00011110110101100011: color_data = 12'b111100000000;
20'b00011110110101100100: color_data = 12'b111100000000;
20'b00011110110101100101: color_data = 12'b111100000000;
20'b00011110110101111101: color_data = 12'b111011101110;
20'b00011110110101111110: color_data = 12'b111011101110;
20'b00011110110101111111: color_data = 12'b111011101110;
20'b00011110110110000000: color_data = 12'b111011101110;
20'b00011110110110000001: color_data = 12'b111011101110;
20'b00011110110110000010: color_data = 12'b111011101110;
20'b00011110110110000011: color_data = 12'b111011101110;
20'b00011110110110000100: color_data = 12'b111011101110;
20'b00011110110110000101: color_data = 12'b111011101110;
20'b00011110110110000110: color_data = 12'b111011101110;
20'b00011110110110001000: color_data = 12'b111011101110;
20'b00011110110110001001: color_data = 12'b111011101110;
20'b00011110110110001010: color_data = 12'b111011101110;
20'b00011110110110001011: color_data = 12'b111011101110;
20'b00011110110110001100: color_data = 12'b111011101110;
20'b00011110110110001101: color_data = 12'b111011101110;
20'b00011110110110001110: color_data = 12'b111011101110;
20'b00011110110110001111: color_data = 12'b111011101110;
20'b00011110110110010000: color_data = 12'b111011101110;
20'b00011110110110010001: color_data = 12'b111011101110;
20'b00011110110110110100: color_data = 12'b111011101110;
20'b00011110110110110101: color_data = 12'b111011101110;
20'b00011110110110110110: color_data = 12'b111011101110;
20'b00011110110110110111: color_data = 12'b111011101110;
20'b00011110110110111000: color_data = 12'b111011101110;
20'b00011110110110111001: color_data = 12'b111011101110;
20'b00011110110110111010: color_data = 12'b111011101110;
20'b00011110110110111011: color_data = 12'b111011101110;
20'b00011110110110111100: color_data = 12'b111011101110;
20'b00011110110110111101: color_data = 12'b111011101110;
20'b00011110110110111111: color_data = 12'b111011101110;
20'b00011110110111000000: color_data = 12'b111011101110;
20'b00011110110111000001: color_data = 12'b111011101110;
20'b00011110110111000010: color_data = 12'b111011101110;
20'b00011110110111000011: color_data = 12'b111011101110;
20'b00011110110111000100: color_data = 12'b111011101110;
20'b00011110110111000101: color_data = 12'b111011101110;
20'b00011110110111000110: color_data = 12'b111011101110;
20'b00011110110111000111: color_data = 12'b111011101110;
20'b00011110110111001000: color_data = 12'b111011101110;
20'b00011110110111001010: color_data = 12'b111011101110;
20'b00011110110111001011: color_data = 12'b111011101110;
20'b00011110110111001100: color_data = 12'b111011101110;
20'b00011110110111001101: color_data = 12'b111011101110;
20'b00011110110111001110: color_data = 12'b111011101110;
20'b00011110110111001111: color_data = 12'b111011101110;
20'b00011110110111010000: color_data = 12'b111011101110;
20'b00011110110111010001: color_data = 12'b111011101110;
20'b00011110110111010010: color_data = 12'b111011101110;
20'b00011110110111010011: color_data = 12'b111011101110;
20'b00011110110111010101: color_data = 12'b111011101110;
20'b00011110110111010110: color_data = 12'b111011101110;
20'b00011110110111010111: color_data = 12'b111011101110;
20'b00011110110111011000: color_data = 12'b111011101110;
20'b00011110110111011001: color_data = 12'b111011101110;
20'b00011110110111011010: color_data = 12'b111011101110;
20'b00011110110111011011: color_data = 12'b111011101110;
20'b00011110110111011100: color_data = 12'b111011101110;
20'b00011110110111011101: color_data = 12'b111011101110;
20'b00011110110111011110: color_data = 12'b111011101110;
20'b00011110110111100000: color_data = 12'b111011101110;
20'b00011110110111100001: color_data = 12'b111011101110;
20'b00011110110111100010: color_data = 12'b111011101110;
20'b00011110110111100011: color_data = 12'b111011101110;
20'b00011110110111100100: color_data = 12'b111011101110;
20'b00011110110111100101: color_data = 12'b111011101110;
20'b00011110110111100110: color_data = 12'b111011101110;
20'b00011110110111100111: color_data = 12'b111011101110;
20'b00011110110111101000: color_data = 12'b111011101110;
20'b00011110110111101001: color_data = 12'b111011101110;
20'b00011111000010101100: color_data = 12'b111011101110;
20'b00011111000010101101: color_data = 12'b111011101110;
20'b00011111000010101110: color_data = 12'b111011101110;
20'b00011111000010101111: color_data = 12'b111011101110;
20'b00011111000010110000: color_data = 12'b111011101110;
20'b00011111000010110001: color_data = 12'b111011101110;
20'b00011111000010110010: color_data = 12'b111011101110;
20'b00011111000010110011: color_data = 12'b111011101110;
20'b00011111000010110100: color_data = 12'b111011101110;
20'b00011111000010110101: color_data = 12'b111011101110;
20'b00011111000010110111: color_data = 12'b111011101110;
20'b00011111000010111000: color_data = 12'b111011101110;
20'b00011111000010111001: color_data = 12'b111011101110;
20'b00011111000010111010: color_data = 12'b111011101110;
20'b00011111000010111011: color_data = 12'b111011101110;
20'b00011111000010111100: color_data = 12'b111011101110;
20'b00011111000010111101: color_data = 12'b111011101110;
20'b00011111000010111110: color_data = 12'b111011101110;
20'b00011111000010111111: color_data = 12'b111011101110;
20'b00011111000011000000: color_data = 12'b111011101110;
20'b00011111000011000010: color_data = 12'b111011101110;
20'b00011111000011000011: color_data = 12'b111011101110;
20'b00011111000011000100: color_data = 12'b111011101110;
20'b00011111000011000101: color_data = 12'b111011101110;
20'b00011111000011000110: color_data = 12'b111011101110;
20'b00011111000011000111: color_data = 12'b111011101110;
20'b00011111000011001000: color_data = 12'b111011101110;
20'b00011111000011001001: color_data = 12'b111011101110;
20'b00011111000011001010: color_data = 12'b111011101110;
20'b00011111000011001011: color_data = 12'b111011101110;
20'b00011111000011001101: color_data = 12'b111011101110;
20'b00011111000011001110: color_data = 12'b111011101110;
20'b00011111000011001111: color_data = 12'b111011101110;
20'b00011111000011010000: color_data = 12'b111011101110;
20'b00011111000011010001: color_data = 12'b111011101110;
20'b00011111000011010010: color_data = 12'b111011101110;
20'b00011111000011010011: color_data = 12'b111011101110;
20'b00011111000011010100: color_data = 12'b111011101110;
20'b00011111000011010101: color_data = 12'b111011101110;
20'b00011111000011010110: color_data = 12'b111011101110;
20'b00011111000100000100: color_data = 12'b111011101110;
20'b00011111000100000101: color_data = 12'b111011101110;
20'b00011111000100000110: color_data = 12'b111011101110;
20'b00011111000100000111: color_data = 12'b111011101110;
20'b00011111000100001000: color_data = 12'b111011101110;
20'b00011111000100001001: color_data = 12'b111011101110;
20'b00011111000100001010: color_data = 12'b111011101110;
20'b00011111000100001011: color_data = 12'b111011101110;
20'b00011111000100001100: color_data = 12'b111011101110;
20'b00011111000100001101: color_data = 12'b111011101110;
20'b00011111000101010001: color_data = 12'b111100000000;
20'b00011111000101010010: color_data = 12'b111100000000;
20'b00011111000101010011: color_data = 12'b111100000000;
20'b00011111000101010100: color_data = 12'b111100000000;
20'b00011111000101010101: color_data = 12'b111100000000;
20'b00011111000101010110: color_data = 12'b111100000000;
20'b00011111000101010111: color_data = 12'b111100000000;
20'b00011111000101011000: color_data = 12'b111100000000;
20'b00011111000101011001: color_data = 12'b111100000000;
20'b00011111000101011010: color_data = 12'b111100000000;
20'b00011111000101011100: color_data = 12'b111100000000;
20'b00011111000101011101: color_data = 12'b111100000000;
20'b00011111000101011110: color_data = 12'b111100000000;
20'b00011111000101011111: color_data = 12'b111100000000;
20'b00011111000101100000: color_data = 12'b111100000000;
20'b00011111000101100001: color_data = 12'b111100000000;
20'b00011111000101100010: color_data = 12'b111100000000;
20'b00011111000101100011: color_data = 12'b111100000000;
20'b00011111000101100100: color_data = 12'b111100000000;
20'b00011111000101100101: color_data = 12'b111100000000;
20'b00011111000101111101: color_data = 12'b111011101110;
20'b00011111000101111110: color_data = 12'b111011101110;
20'b00011111000101111111: color_data = 12'b111011101110;
20'b00011111000110000000: color_data = 12'b111011101110;
20'b00011111000110000001: color_data = 12'b111011101110;
20'b00011111000110000010: color_data = 12'b111011101110;
20'b00011111000110000011: color_data = 12'b111011101110;
20'b00011111000110000100: color_data = 12'b111011101110;
20'b00011111000110000101: color_data = 12'b111011101110;
20'b00011111000110000110: color_data = 12'b111011101110;
20'b00011111000110001000: color_data = 12'b111011101110;
20'b00011111000110001001: color_data = 12'b111011101110;
20'b00011111000110001010: color_data = 12'b111011101110;
20'b00011111000110001011: color_data = 12'b111011101110;
20'b00011111000110001100: color_data = 12'b111011101110;
20'b00011111000110001101: color_data = 12'b111011101110;
20'b00011111000110001110: color_data = 12'b111011101110;
20'b00011111000110001111: color_data = 12'b111011101110;
20'b00011111000110010000: color_data = 12'b111011101110;
20'b00011111000110010001: color_data = 12'b111011101110;
20'b00011111000110110100: color_data = 12'b111011101110;
20'b00011111000110110101: color_data = 12'b111011101110;
20'b00011111000110110110: color_data = 12'b111011101110;
20'b00011111000110110111: color_data = 12'b111011101110;
20'b00011111000110111000: color_data = 12'b111011101110;
20'b00011111000110111001: color_data = 12'b111011101110;
20'b00011111000110111010: color_data = 12'b111011101110;
20'b00011111000110111011: color_data = 12'b111011101110;
20'b00011111000110111100: color_data = 12'b111011101110;
20'b00011111000110111101: color_data = 12'b111011101110;
20'b00011111000110111111: color_data = 12'b111011101110;
20'b00011111000111000000: color_data = 12'b111011101110;
20'b00011111000111000001: color_data = 12'b111011101110;
20'b00011111000111000010: color_data = 12'b111011101110;
20'b00011111000111000011: color_data = 12'b111011101110;
20'b00011111000111000100: color_data = 12'b111011101110;
20'b00011111000111000101: color_data = 12'b111011101110;
20'b00011111000111000110: color_data = 12'b111011101110;
20'b00011111000111000111: color_data = 12'b111011101110;
20'b00011111000111001000: color_data = 12'b111011101110;
20'b00011111000111001010: color_data = 12'b111011101110;
20'b00011111000111001011: color_data = 12'b111011101110;
20'b00011111000111001100: color_data = 12'b111011101110;
20'b00011111000111001101: color_data = 12'b111011101110;
20'b00011111000111001110: color_data = 12'b111011101110;
20'b00011111000111001111: color_data = 12'b111011101110;
20'b00011111000111010000: color_data = 12'b111011101110;
20'b00011111000111010001: color_data = 12'b111011101110;
20'b00011111000111010010: color_data = 12'b111011101110;
20'b00011111000111010011: color_data = 12'b111011101110;
20'b00011111000111010101: color_data = 12'b111011101110;
20'b00011111000111010110: color_data = 12'b111011101110;
20'b00011111000111010111: color_data = 12'b111011101110;
20'b00011111000111011000: color_data = 12'b111011101110;
20'b00011111000111011001: color_data = 12'b111011101110;
20'b00011111000111011010: color_data = 12'b111011101110;
20'b00011111000111011011: color_data = 12'b111011101110;
20'b00011111000111011100: color_data = 12'b111011101110;
20'b00011111000111011101: color_data = 12'b111011101110;
20'b00011111000111011110: color_data = 12'b111011101110;
20'b00011111000111100000: color_data = 12'b111011101110;
20'b00011111000111100001: color_data = 12'b111011101110;
20'b00011111000111100010: color_data = 12'b111011101110;
20'b00011111000111100011: color_data = 12'b111011101110;
20'b00011111000111100100: color_data = 12'b111011101110;
20'b00011111000111100101: color_data = 12'b111011101110;
20'b00011111000111100110: color_data = 12'b111011101110;
20'b00011111000111100111: color_data = 12'b111011101110;
20'b00011111000111101000: color_data = 12'b111011101110;
20'b00011111000111101001: color_data = 12'b111011101110;
20'b00011111010110110100: color_data = 12'b111011101110;
20'b00011111010110110101: color_data = 12'b111011101110;
20'b00011111010110110110: color_data = 12'b111011101110;
20'b00011111010110110111: color_data = 12'b111011101110;
20'b00011111010110111000: color_data = 12'b111011101110;
20'b00011111010110111001: color_data = 12'b111011101110;
20'b00011111010110111010: color_data = 12'b111011101110;
20'b00011111010110111011: color_data = 12'b111011101110;
20'b00011111010110111100: color_data = 12'b111011101110;
20'b00011111010110111101: color_data = 12'b111011101110;
20'b00011111010110111111: color_data = 12'b111011101110;
20'b00011111010111000000: color_data = 12'b111011101110;
20'b00011111010111000001: color_data = 12'b111011101110;
20'b00011111010111000010: color_data = 12'b111011101110;
20'b00011111010111000011: color_data = 12'b111011101110;
20'b00011111010111000100: color_data = 12'b111011101110;
20'b00011111010111000101: color_data = 12'b111011101110;
20'b00011111010111000110: color_data = 12'b111011101110;
20'b00011111010111000111: color_data = 12'b111011101110;
20'b00011111010111001000: color_data = 12'b111011101110;
20'b00011111010111001010: color_data = 12'b111011101110;
20'b00011111010111001011: color_data = 12'b111011101110;
20'b00011111010111001100: color_data = 12'b111011101110;
20'b00011111010111001101: color_data = 12'b111011101110;
20'b00011111010111001110: color_data = 12'b111011101110;
20'b00011111010111001111: color_data = 12'b111011101110;
20'b00011111010111010000: color_data = 12'b111011101110;
20'b00011111010111010001: color_data = 12'b111011101110;
20'b00011111010111010010: color_data = 12'b111011101110;
20'b00011111010111010011: color_data = 12'b111011101110;
20'b00011111010111010101: color_data = 12'b111011101110;
20'b00011111010111010110: color_data = 12'b111011101110;
20'b00011111010111010111: color_data = 12'b111011101110;
20'b00011111010111011000: color_data = 12'b111011101110;
20'b00011111010111011001: color_data = 12'b111011101110;
20'b00011111010111011010: color_data = 12'b111011101110;
20'b00011111010111011011: color_data = 12'b111011101110;
20'b00011111010111011100: color_data = 12'b111011101110;
20'b00011111010111011101: color_data = 12'b111011101110;
20'b00011111010111011110: color_data = 12'b111011101110;
20'b00011111010111100000: color_data = 12'b111011101110;
20'b00011111010111100001: color_data = 12'b111011101110;
20'b00011111010111100010: color_data = 12'b111011101110;
20'b00011111010111100011: color_data = 12'b111011101110;
20'b00011111010111100100: color_data = 12'b111011101110;
20'b00011111010111100101: color_data = 12'b111011101110;
20'b00011111010111100110: color_data = 12'b111011101110;
20'b00011111010111100111: color_data = 12'b111011101110;
20'b00011111010111101000: color_data = 12'b111011101110;
20'b00011111010111101001: color_data = 12'b111011101110;
20'b00011111100011001101: color_data = 12'b111011101110;
20'b00011111100011001110: color_data = 12'b111011101110;
20'b00011111100011001111: color_data = 12'b111011101110;
20'b00011111100011010000: color_data = 12'b111011101110;
20'b00011111100011010001: color_data = 12'b111011101110;
20'b00011111100011010010: color_data = 12'b111011101110;
20'b00011111100011010011: color_data = 12'b111011101110;
20'b00011111100011010100: color_data = 12'b111011101110;
20'b00011111100011010101: color_data = 12'b111011101110;
20'b00011111100011010110: color_data = 12'b111011101110;
20'b00011111100011011000: color_data = 12'b111011101110;
20'b00011111100011011001: color_data = 12'b111011101110;
20'b00011111100011011010: color_data = 12'b111011101110;
20'b00011111100011011011: color_data = 12'b111011101110;
20'b00011111100011011100: color_data = 12'b111011101110;
20'b00011111100011011101: color_data = 12'b111011101110;
20'b00011111100011011110: color_data = 12'b111011101110;
20'b00011111100011011111: color_data = 12'b111011101110;
20'b00011111100011100000: color_data = 12'b111011101110;
20'b00011111100011100001: color_data = 12'b111011101110;
20'b00011111100011111001: color_data = 12'b111011101110;
20'b00011111100011111010: color_data = 12'b111011101110;
20'b00011111100011111011: color_data = 12'b111011101110;
20'b00011111100011111100: color_data = 12'b111011101110;
20'b00011111100011111101: color_data = 12'b111011101110;
20'b00011111100011111110: color_data = 12'b111011101110;
20'b00011111100011111111: color_data = 12'b111011101110;
20'b00011111100100000000: color_data = 12'b111011101110;
20'b00011111100100000001: color_data = 12'b111011101110;
20'b00011111100100000010: color_data = 12'b111011101110;
20'b00011111100100000100: color_data = 12'b111011101110;
20'b00011111100100000101: color_data = 12'b111011101110;
20'b00011111100100000110: color_data = 12'b111011101110;
20'b00011111100100000111: color_data = 12'b111011101110;
20'b00011111100100001000: color_data = 12'b111011101110;
20'b00011111100100001001: color_data = 12'b111011101110;
20'b00011111100100001010: color_data = 12'b111011101110;
20'b00011111100100001011: color_data = 12'b111011101110;
20'b00011111100100001100: color_data = 12'b111011101110;
20'b00011111100100001101: color_data = 12'b111011101110;
20'b00011111100100100101: color_data = 12'b111011101110;
20'b00011111100100100110: color_data = 12'b111011101110;
20'b00011111100100100111: color_data = 12'b111011101110;
20'b00011111100100101000: color_data = 12'b111011101110;
20'b00011111100100101001: color_data = 12'b111011101110;
20'b00011111100100101010: color_data = 12'b111011101110;
20'b00011111100100101011: color_data = 12'b111011101110;
20'b00011111100100101100: color_data = 12'b111011101110;
20'b00011111100100101101: color_data = 12'b111011101110;
20'b00011111100100101110: color_data = 12'b111011101110;
20'b00011111100101000110: color_data = 12'b111011101110;
20'b00011111100101000111: color_data = 12'b111011101110;
20'b00011111100101001000: color_data = 12'b111011101110;
20'b00011111100101001001: color_data = 12'b111011101110;
20'b00011111100101001010: color_data = 12'b111011101110;
20'b00011111100101001011: color_data = 12'b111011101110;
20'b00011111100101001100: color_data = 12'b111011101110;
20'b00011111100101001101: color_data = 12'b111011101110;
20'b00011111100101001110: color_data = 12'b111011101110;
20'b00011111100101001111: color_data = 12'b111011101110;
20'b00011111100101110010: color_data = 12'b111011101110;
20'b00011111100101110011: color_data = 12'b111011101110;
20'b00011111100101110100: color_data = 12'b111011101110;
20'b00011111100101110101: color_data = 12'b111011101110;
20'b00011111100101110110: color_data = 12'b111011101110;
20'b00011111100101110111: color_data = 12'b111011101110;
20'b00011111100101111000: color_data = 12'b111011101110;
20'b00011111100101111001: color_data = 12'b111011101110;
20'b00011111100101111010: color_data = 12'b111011101110;
20'b00011111100101111011: color_data = 12'b111011101110;
20'b00011111100101111101: color_data = 12'b111011101110;
20'b00011111100101111110: color_data = 12'b111011101110;
20'b00011111100101111111: color_data = 12'b111011101110;
20'b00011111100110000000: color_data = 12'b111011101110;
20'b00011111100110000001: color_data = 12'b111011101110;
20'b00011111100110000010: color_data = 12'b111011101110;
20'b00011111100110000011: color_data = 12'b111011101110;
20'b00011111100110000100: color_data = 12'b111011101110;
20'b00011111100110000101: color_data = 12'b111011101110;
20'b00011111100110000110: color_data = 12'b111011101110;
20'b00011111100110001000: color_data = 12'b111011101110;
20'b00011111100110001001: color_data = 12'b111011101110;
20'b00011111100110001010: color_data = 12'b111011101110;
20'b00011111100110001011: color_data = 12'b111011101110;
20'b00011111100110001100: color_data = 12'b111011101110;
20'b00011111100110001101: color_data = 12'b111011101110;
20'b00011111100110001110: color_data = 12'b111011101110;
20'b00011111100110001111: color_data = 12'b111011101110;
20'b00011111100110010000: color_data = 12'b111011101110;
20'b00011111100110010001: color_data = 12'b111011101110;
20'b00011111110011001101: color_data = 12'b111011101110;
20'b00011111110011001110: color_data = 12'b111011101110;
20'b00011111110011001111: color_data = 12'b111011101110;
20'b00011111110011010000: color_data = 12'b111011101110;
20'b00011111110011010001: color_data = 12'b111011101110;
20'b00011111110011010010: color_data = 12'b111011101110;
20'b00011111110011010011: color_data = 12'b111011101110;
20'b00011111110011010100: color_data = 12'b111011101110;
20'b00011111110011010101: color_data = 12'b111011101110;
20'b00011111110011010110: color_data = 12'b111011101110;
20'b00011111110011011000: color_data = 12'b111011101110;
20'b00011111110011011001: color_data = 12'b111011101110;
20'b00011111110011011010: color_data = 12'b111011101110;
20'b00011111110011011011: color_data = 12'b111011101110;
20'b00011111110011011100: color_data = 12'b111011101110;
20'b00011111110011011101: color_data = 12'b111011101110;
20'b00011111110011011110: color_data = 12'b111011101110;
20'b00011111110011011111: color_data = 12'b111011101110;
20'b00011111110011100000: color_data = 12'b111011101110;
20'b00011111110011100001: color_data = 12'b111011101110;
20'b00011111110011111001: color_data = 12'b111011101110;
20'b00011111110011111010: color_data = 12'b111011101110;
20'b00011111110011111011: color_data = 12'b111011101110;
20'b00011111110011111100: color_data = 12'b111011101110;
20'b00011111110011111101: color_data = 12'b111011101110;
20'b00011111110011111110: color_data = 12'b111011101110;
20'b00011111110011111111: color_data = 12'b111011101110;
20'b00011111110100000000: color_data = 12'b111011101110;
20'b00011111110100000001: color_data = 12'b111011101110;
20'b00011111110100000010: color_data = 12'b111011101110;
20'b00011111110100000100: color_data = 12'b111011101110;
20'b00011111110100000101: color_data = 12'b111011101110;
20'b00011111110100000110: color_data = 12'b111011101110;
20'b00011111110100000111: color_data = 12'b111011101110;
20'b00011111110100001000: color_data = 12'b111011101110;
20'b00011111110100001001: color_data = 12'b111011101110;
20'b00011111110100001010: color_data = 12'b111011101110;
20'b00011111110100001011: color_data = 12'b111011101110;
20'b00011111110100001100: color_data = 12'b111011101110;
20'b00011111110100001101: color_data = 12'b111011101110;
20'b00011111110100100101: color_data = 12'b111011101110;
20'b00011111110100100110: color_data = 12'b111011101110;
20'b00011111110100100111: color_data = 12'b111011101110;
20'b00011111110100101000: color_data = 12'b111011101110;
20'b00011111110100101001: color_data = 12'b111011101110;
20'b00011111110100101010: color_data = 12'b111011101110;
20'b00011111110100101011: color_data = 12'b111011101110;
20'b00011111110100101100: color_data = 12'b111011101110;
20'b00011111110100101101: color_data = 12'b111011101110;
20'b00011111110100101110: color_data = 12'b111011101110;
20'b00011111110101000110: color_data = 12'b111011101110;
20'b00011111110101000111: color_data = 12'b111011101110;
20'b00011111110101001000: color_data = 12'b111011101110;
20'b00011111110101001001: color_data = 12'b111011101110;
20'b00011111110101001010: color_data = 12'b111011101110;
20'b00011111110101001011: color_data = 12'b111011101110;
20'b00011111110101001100: color_data = 12'b111011101110;
20'b00011111110101001101: color_data = 12'b111011101110;
20'b00011111110101001110: color_data = 12'b111011101110;
20'b00011111110101001111: color_data = 12'b111011101110;
20'b00011111110101110010: color_data = 12'b111011101110;
20'b00011111110101110011: color_data = 12'b111011101110;
20'b00011111110101110100: color_data = 12'b111011101110;
20'b00011111110101110101: color_data = 12'b111011101110;
20'b00011111110101110110: color_data = 12'b111011101110;
20'b00011111110101110111: color_data = 12'b111011101110;
20'b00011111110101111000: color_data = 12'b111011101110;
20'b00011111110101111001: color_data = 12'b111011101110;
20'b00011111110101111010: color_data = 12'b111011101110;
20'b00011111110101111011: color_data = 12'b111011101110;
20'b00011111110101111101: color_data = 12'b111011101110;
20'b00011111110101111110: color_data = 12'b111011101110;
20'b00011111110101111111: color_data = 12'b111011101110;
20'b00011111110110000000: color_data = 12'b111011101110;
20'b00011111110110000001: color_data = 12'b111011101110;
20'b00011111110110000010: color_data = 12'b111011101110;
20'b00011111110110000011: color_data = 12'b111011101110;
20'b00011111110110000100: color_data = 12'b111011101110;
20'b00011111110110000101: color_data = 12'b111011101110;
20'b00011111110110000110: color_data = 12'b111011101110;
20'b00011111110110001000: color_data = 12'b111011101110;
20'b00011111110110001001: color_data = 12'b111011101110;
20'b00011111110110001010: color_data = 12'b111011101110;
20'b00011111110110001011: color_data = 12'b111011101110;
20'b00011111110110001100: color_data = 12'b111011101110;
20'b00011111110110001101: color_data = 12'b111011101110;
20'b00011111110110001110: color_data = 12'b111011101110;
20'b00011111110110001111: color_data = 12'b111011101110;
20'b00011111110110010000: color_data = 12'b111011101110;
20'b00011111110110010001: color_data = 12'b111011101110;
20'b00011111110110101001: color_data = 12'b111011101110;
20'b00011111110110101010: color_data = 12'b111011101110;
20'b00011111110110101011: color_data = 12'b111011101110;
20'b00011111110110101100: color_data = 12'b111011101110;
20'b00011111110110101101: color_data = 12'b111011101110;
20'b00011111110110101110: color_data = 12'b111011101110;
20'b00011111110110101111: color_data = 12'b111011101110;
20'b00011111110110110000: color_data = 12'b111011101110;
20'b00011111110110110001: color_data = 12'b111011101110;
20'b00011111110110110010: color_data = 12'b111011101110;
20'b00100000000011001101: color_data = 12'b111011101110;
20'b00100000000011001110: color_data = 12'b111011101110;
20'b00100000000011001111: color_data = 12'b111011101110;
20'b00100000000011010000: color_data = 12'b111011101110;
20'b00100000000011010001: color_data = 12'b111011101110;
20'b00100000000011010010: color_data = 12'b111011101110;
20'b00100000000011010011: color_data = 12'b111011101110;
20'b00100000000011010100: color_data = 12'b111011101110;
20'b00100000000011010101: color_data = 12'b111011101110;
20'b00100000000011010110: color_data = 12'b111011101110;
20'b00100000000011011000: color_data = 12'b111011101110;
20'b00100000000011011001: color_data = 12'b111011101110;
20'b00100000000011011010: color_data = 12'b111011101110;
20'b00100000000011011011: color_data = 12'b111011101110;
20'b00100000000011011100: color_data = 12'b111011101110;
20'b00100000000011011101: color_data = 12'b111011101110;
20'b00100000000011011110: color_data = 12'b111011101110;
20'b00100000000011011111: color_data = 12'b111011101110;
20'b00100000000011100000: color_data = 12'b111011101110;
20'b00100000000011100001: color_data = 12'b111011101110;
20'b00100000000011111001: color_data = 12'b111011101110;
20'b00100000000011111010: color_data = 12'b111011101110;
20'b00100000000011111011: color_data = 12'b111011101110;
20'b00100000000011111100: color_data = 12'b111011101110;
20'b00100000000011111101: color_data = 12'b111011101110;
20'b00100000000011111110: color_data = 12'b111011101110;
20'b00100000000011111111: color_data = 12'b111011101110;
20'b00100000000100000000: color_data = 12'b111011101110;
20'b00100000000100000001: color_data = 12'b111011101110;
20'b00100000000100000010: color_data = 12'b111011101110;
20'b00100000000100000100: color_data = 12'b111011101110;
20'b00100000000100000101: color_data = 12'b111011101110;
20'b00100000000100000110: color_data = 12'b111011101110;
20'b00100000000100000111: color_data = 12'b111011101110;
20'b00100000000100001000: color_data = 12'b111011101110;
20'b00100000000100001001: color_data = 12'b111011101110;
20'b00100000000100001010: color_data = 12'b111011101110;
20'b00100000000100001011: color_data = 12'b111011101110;
20'b00100000000100001100: color_data = 12'b111011101110;
20'b00100000000100001101: color_data = 12'b111011101110;
20'b00100000000100100101: color_data = 12'b111011101110;
20'b00100000000100100110: color_data = 12'b111011101110;
20'b00100000000100100111: color_data = 12'b111011101110;
20'b00100000000100101000: color_data = 12'b111011101110;
20'b00100000000100101001: color_data = 12'b111011101110;
20'b00100000000100101010: color_data = 12'b111011101110;
20'b00100000000100101011: color_data = 12'b111011101110;
20'b00100000000100101100: color_data = 12'b111011101110;
20'b00100000000100101101: color_data = 12'b111011101110;
20'b00100000000100101110: color_data = 12'b111011101110;
20'b00100000000101000110: color_data = 12'b111011101110;
20'b00100000000101000111: color_data = 12'b111011101110;
20'b00100000000101001000: color_data = 12'b111011101110;
20'b00100000000101001001: color_data = 12'b111011101110;
20'b00100000000101001010: color_data = 12'b111011101110;
20'b00100000000101001011: color_data = 12'b111011101110;
20'b00100000000101001100: color_data = 12'b111011101110;
20'b00100000000101001101: color_data = 12'b111011101110;
20'b00100000000101001110: color_data = 12'b111011101110;
20'b00100000000101001111: color_data = 12'b111011101110;
20'b00100000000101110010: color_data = 12'b111011101110;
20'b00100000000101110011: color_data = 12'b111011101110;
20'b00100000000101110100: color_data = 12'b111011101110;
20'b00100000000101110101: color_data = 12'b111011101110;
20'b00100000000101110110: color_data = 12'b111011101110;
20'b00100000000101110111: color_data = 12'b111011101110;
20'b00100000000101111000: color_data = 12'b111011101110;
20'b00100000000101111001: color_data = 12'b111011101110;
20'b00100000000101111010: color_data = 12'b111011101110;
20'b00100000000101111011: color_data = 12'b111011101110;
20'b00100000000101111101: color_data = 12'b111011101110;
20'b00100000000101111110: color_data = 12'b111011101110;
20'b00100000000101111111: color_data = 12'b111011101110;
20'b00100000000110000000: color_data = 12'b111011101110;
20'b00100000000110000001: color_data = 12'b111011101110;
20'b00100000000110000010: color_data = 12'b111011101110;
20'b00100000000110000011: color_data = 12'b111011101110;
20'b00100000000110000100: color_data = 12'b111011101110;
20'b00100000000110000101: color_data = 12'b111011101110;
20'b00100000000110000110: color_data = 12'b111011101110;
20'b00100000000110001000: color_data = 12'b111011101110;
20'b00100000000110001001: color_data = 12'b111011101110;
20'b00100000000110001010: color_data = 12'b111011101110;
20'b00100000000110001011: color_data = 12'b111011101110;
20'b00100000000110001100: color_data = 12'b111011101110;
20'b00100000000110001101: color_data = 12'b111011101110;
20'b00100000000110001110: color_data = 12'b111011101110;
20'b00100000000110001111: color_data = 12'b111011101110;
20'b00100000000110010000: color_data = 12'b111011101110;
20'b00100000000110010001: color_data = 12'b111011101110;
20'b00100000000110101001: color_data = 12'b111011101110;
20'b00100000000110101010: color_data = 12'b111011101110;
20'b00100000000110101011: color_data = 12'b111011101110;
20'b00100000000110101100: color_data = 12'b111011101110;
20'b00100000000110101101: color_data = 12'b111011101110;
20'b00100000000110101110: color_data = 12'b111011101110;
20'b00100000000110101111: color_data = 12'b111011101110;
20'b00100000000110110000: color_data = 12'b111011101110;
20'b00100000000110110001: color_data = 12'b111011101110;
20'b00100000000110110010: color_data = 12'b111011101110;
20'b00100000010011001101: color_data = 12'b111011101110;
20'b00100000010011001110: color_data = 12'b111011101110;
20'b00100000010011001111: color_data = 12'b111011101110;
20'b00100000010011010000: color_data = 12'b111011101110;
20'b00100000010011010001: color_data = 12'b111011101110;
20'b00100000010011010010: color_data = 12'b111011101110;
20'b00100000010011010011: color_data = 12'b111011101110;
20'b00100000010011010100: color_data = 12'b111011101110;
20'b00100000010011010101: color_data = 12'b111011101110;
20'b00100000010011010110: color_data = 12'b111011101110;
20'b00100000010011011000: color_data = 12'b111011101110;
20'b00100000010011011001: color_data = 12'b111011101110;
20'b00100000010011011010: color_data = 12'b111011101110;
20'b00100000010011011011: color_data = 12'b111011101110;
20'b00100000010011011100: color_data = 12'b111011101110;
20'b00100000010011011101: color_data = 12'b111011101110;
20'b00100000010011011110: color_data = 12'b111011101110;
20'b00100000010011011111: color_data = 12'b111011101110;
20'b00100000010011100000: color_data = 12'b111011101110;
20'b00100000010011100001: color_data = 12'b111011101110;
20'b00100000010011111001: color_data = 12'b111011101110;
20'b00100000010011111010: color_data = 12'b111011101110;
20'b00100000010011111011: color_data = 12'b111011101110;
20'b00100000010011111100: color_data = 12'b111011101110;
20'b00100000010011111101: color_data = 12'b111011101110;
20'b00100000010011111110: color_data = 12'b111011101110;
20'b00100000010011111111: color_data = 12'b111011101110;
20'b00100000010100000000: color_data = 12'b111011101110;
20'b00100000010100000001: color_data = 12'b111011101110;
20'b00100000010100000010: color_data = 12'b111011101110;
20'b00100000010100000100: color_data = 12'b111011101110;
20'b00100000010100000101: color_data = 12'b111011101110;
20'b00100000010100000110: color_data = 12'b111011101110;
20'b00100000010100000111: color_data = 12'b111011101110;
20'b00100000010100001000: color_data = 12'b111011101110;
20'b00100000010100001001: color_data = 12'b111011101110;
20'b00100000010100001010: color_data = 12'b111011101110;
20'b00100000010100001011: color_data = 12'b111011101110;
20'b00100000010100001100: color_data = 12'b111011101110;
20'b00100000010100001101: color_data = 12'b111011101110;
20'b00100000010100100101: color_data = 12'b111011101110;
20'b00100000010100100110: color_data = 12'b111011101110;
20'b00100000010100100111: color_data = 12'b111011101110;
20'b00100000010100101000: color_data = 12'b111011101110;
20'b00100000010100101001: color_data = 12'b111011101110;
20'b00100000010100101010: color_data = 12'b111011101110;
20'b00100000010100101011: color_data = 12'b111011101110;
20'b00100000010100101100: color_data = 12'b111011101110;
20'b00100000010100101101: color_data = 12'b111011101110;
20'b00100000010100101110: color_data = 12'b111011101110;
20'b00100000010101000110: color_data = 12'b111011101110;
20'b00100000010101000111: color_data = 12'b111011101110;
20'b00100000010101001000: color_data = 12'b111011101110;
20'b00100000010101001001: color_data = 12'b111011101110;
20'b00100000010101001010: color_data = 12'b111011101110;
20'b00100000010101001011: color_data = 12'b111011101110;
20'b00100000010101001100: color_data = 12'b111011101110;
20'b00100000010101001101: color_data = 12'b111011101110;
20'b00100000010101001110: color_data = 12'b111011101110;
20'b00100000010101001111: color_data = 12'b111011101110;
20'b00100000010101110010: color_data = 12'b111011101110;
20'b00100000010101110011: color_data = 12'b111011101110;
20'b00100000010101110100: color_data = 12'b111011101110;
20'b00100000010101110101: color_data = 12'b111011101110;
20'b00100000010101110110: color_data = 12'b111011101110;
20'b00100000010101110111: color_data = 12'b111011101110;
20'b00100000010101111000: color_data = 12'b111011101110;
20'b00100000010101111001: color_data = 12'b111011101110;
20'b00100000010101111010: color_data = 12'b111011101110;
20'b00100000010101111011: color_data = 12'b111011101110;
20'b00100000010101111101: color_data = 12'b111011101110;
20'b00100000010101111110: color_data = 12'b111011101110;
20'b00100000010101111111: color_data = 12'b111011101110;
20'b00100000010110000000: color_data = 12'b111011101110;
20'b00100000010110000001: color_data = 12'b111011101110;
20'b00100000010110000010: color_data = 12'b111011101110;
20'b00100000010110000011: color_data = 12'b111011101110;
20'b00100000010110000100: color_data = 12'b111011101110;
20'b00100000010110000101: color_data = 12'b111011101110;
20'b00100000010110000110: color_data = 12'b111011101110;
20'b00100000010110001000: color_data = 12'b111011101110;
20'b00100000010110001001: color_data = 12'b111011101110;
20'b00100000010110001010: color_data = 12'b111011101110;
20'b00100000010110001011: color_data = 12'b111011101110;
20'b00100000010110001100: color_data = 12'b111011101110;
20'b00100000010110001101: color_data = 12'b111011101110;
20'b00100000010110001110: color_data = 12'b111011101110;
20'b00100000010110001111: color_data = 12'b111011101110;
20'b00100000010110010000: color_data = 12'b111011101110;
20'b00100000010110010001: color_data = 12'b111011101110;
20'b00100000010110101001: color_data = 12'b111011101110;
20'b00100000010110101010: color_data = 12'b111011101110;
20'b00100000010110101011: color_data = 12'b111011101110;
20'b00100000010110101100: color_data = 12'b111011101110;
20'b00100000010110101101: color_data = 12'b111011101110;
20'b00100000010110101110: color_data = 12'b111011101110;
20'b00100000010110101111: color_data = 12'b111011101110;
20'b00100000010110110000: color_data = 12'b111011101110;
20'b00100000010110110001: color_data = 12'b111011101110;
20'b00100000010110110010: color_data = 12'b111011101110;
20'b00100000100011001101: color_data = 12'b111011101110;
20'b00100000100011001110: color_data = 12'b111011101110;
20'b00100000100011001111: color_data = 12'b111011101110;
20'b00100000100011010000: color_data = 12'b111011101110;
20'b00100000100011010001: color_data = 12'b111011101110;
20'b00100000100011010010: color_data = 12'b111011101110;
20'b00100000100011010011: color_data = 12'b111011101110;
20'b00100000100011010100: color_data = 12'b111011101110;
20'b00100000100011010101: color_data = 12'b111011101110;
20'b00100000100011010110: color_data = 12'b111011101110;
20'b00100000100011011000: color_data = 12'b111011101110;
20'b00100000100011011001: color_data = 12'b111011101110;
20'b00100000100011011010: color_data = 12'b111011101110;
20'b00100000100011011011: color_data = 12'b111011101110;
20'b00100000100011011100: color_data = 12'b111011101110;
20'b00100000100011011101: color_data = 12'b111011101110;
20'b00100000100011011110: color_data = 12'b111011101110;
20'b00100000100011011111: color_data = 12'b111011101110;
20'b00100000100011100000: color_data = 12'b111011101110;
20'b00100000100011100001: color_data = 12'b111011101110;
20'b00100000100011111001: color_data = 12'b111011101110;
20'b00100000100011111010: color_data = 12'b111011101110;
20'b00100000100011111011: color_data = 12'b111011101110;
20'b00100000100011111100: color_data = 12'b111011101110;
20'b00100000100011111101: color_data = 12'b111011101110;
20'b00100000100011111110: color_data = 12'b111011101110;
20'b00100000100011111111: color_data = 12'b111011101110;
20'b00100000100100000000: color_data = 12'b111011101110;
20'b00100000100100000001: color_data = 12'b111011101110;
20'b00100000100100000010: color_data = 12'b111011101110;
20'b00100000100100000100: color_data = 12'b111011101110;
20'b00100000100100000101: color_data = 12'b111011101110;
20'b00100000100100000110: color_data = 12'b111011101110;
20'b00100000100100000111: color_data = 12'b111011101110;
20'b00100000100100001000: color_data = 12'b111011101110;
20'b00100000100100001001: color_data = 12'b111011101110;
20'b00100000100100001010: color_data = 12'b111011101110;
20'b00100000100100001011: color_data = 12'b111011101110;
20'b00100000100100001100: color_data = 12'b111011101110;
20'b00100000100100001101: color_data = 12'b111011101110;
20'b00100000100100100101: color_data = 12'b111011101110;
20'b00100000100100100110: color_data = 12'b111011101110;
20'b00100000100100100111: color_data = 12'b111011101110;
20'b00100000100100101000: color_data = 12'b111011101110;
20'b00100000100100101001: color_data = 12'b111011101110;
20'b00100000100100101010: color_data = 12'b111011101110;
20'b00100000100100101011: color_data = 12'b111011101110;
20'b00100000100100101100: color_data = 12'b111011101110;
20'b00100000100100101101: color_data = 12'b111011101110;
20'b00100000100100101110: color_data = 12'b111011101110;
20'b00100000100101000110: color_data = 12'b111011101110;
20'b00100000100101000111: color_data = 12'b111011101110;
20'b00100000100101001000: color_data = 12'b111011101110;
20'b00100000100101001001: color_data = 12'b111011101110;
20'b00100000100101001010: color_data = 12'b111011101110;
20'b00100000100101001011: color_data = 12'b111011101110;
20'b00100000100101001100: color_data = 12'b111011101110;
20'b00100000100101001101: color_data = 12'b111011101110;
20'b00100000100101001110: color_data = 12'b111011101110;
20'b00100000100101001111: color_data = 12'b111011101110;
20'b00100000100101110010: color_data = 12'b111011101110;
20'b00100000100101110011: color_data = 12'b111011101110;
20'b00100000100101110100: color_data = 12'b111011101110;
20'b00100000100101110101: color_data = 12'b111011101110;
20'b00100000100101110110: color_data = 12'b111011101110;
20'b00100000100101110111: color_data = 12'b111011101110;
20'b00100000100101111000: color_data = 12'b111011101110;
20'b00100000100101111001: color_data = 12'b111011101110;
20'b00100000100101111010: color_data = 12'b111011101110;
20'b00100000100101111011: color_data = 12'b111011101110;
20'b00100000100101111101: color_data = 12'b111011101110;
20'b00100000100101111110: color_data = 12'b111011101110;
20'b00100000100101111111: color_data = 12'b111011101110;
20'b00100000100110000000: color_data = 12'b111011101110;
20'b00100000100110000001: color_data = 12'b111011101110;
20'b00100000100110000010: color_data = 12'b111011101110;
20'b00100000100110000011: color_data = 12'b111011101110;
20'b00100000100110000100: color_data = 12'b111011101110;
20'b00100000100110000101: color_data = 12'b111011101110;
20'b00100000100110000110: color_data = 12'b111011101110;
20'b00100000100110001000: color_data = 12'b111011101110;
20'b00100000100110001001: color_data = 12'b111011101110;
20'b00100000100110001010: color_data = 12'b111011101110;
20'b00100000100110001011: color_data = 12'b111011101110;
20'b00100000100110001100: color_data = 12'b111011101110;
20'b00100000100110001101: color_data = 12'b111011101110;
20'b00100000100110001110: color_data = 12'b111011101110;
20'b00100000100110001111: color_data = 12'b111011101110;
20'b00100000100110010000: color_data = 12'b111011101110;
20'b00100000100110010001: color_data = 12'b111011101110;
20'b00100000100110101001: color_data = 12'b111011101110;
20'b00100000100110101010: color_data = 12'b111011101110;
20'b00100000100110101011: color_data = 12'b111011101110;
20'b00100000100110101100: color_data = 12'b111011101110;
20'b00100000100110101101: color_data = 12'b111011101110;
20'b00100000100110101110: color_data = 12'b111011101110;
20'b00100000100110101111: color_data = 12'b111011101110;
20'b00100000100110110000: color_data = 12'b111011101110;
20'b00100000100110110001: color_data = 12'b111011101110;
20'b00100000100110110010: color_data = 12'b111011101110;
20'b00100000110011001101: color_data = 12'b111011101110;
20'b00100000110011001110: color_data = 12'b111011101110;
20'b00100000110011001111: color_data = 12'b111011101110;
20'b00100000110011010000: color_data = 12'b111011101110;
20'b00100000110011010001: color_data = 12'b111011101110;
20'b00100000110011010010: color_data = 12'b111011101110;
20'b00100000110011010011: color_data = 12'b111011101110;
20'b00100000110011010100: color_data = 12'b111011101110;
20'b00100000110011010101: color_data = 12'b111011101110;
20'b00100000110011010110: color_data = 12'b111011101110;
20'b00100000110011011000: color_data = 12'b111011101110;
20'b00100000110011011001: color_data = 12'b111011101110;
20'b00100000110011011010: color_data = 12'b111011101110;
20'b00100000110011011011: color_data = 12'b111011101110;
20'b00100000110011011100: color_data = 12'b111011101110;
20'b00100000110011011101: color_data = 12'b111011101110;
20'b00100000110011011110: color_data = 12'b111011101110;
20'b00100000110011011111: color_data = 12'b111011101110;
20'b00100000110011100000: color_data = 12'b111011101110;
20'b00100000110011100001: color_data = 12'b111011101110;
20'b00100000110011111001: color_data = 12'b111011101110;
20'b00100000110011111010: color_data = 12'b111011101110;
20'b00100000110011111011: color_data = 12'b111011101110;
20'b00100000110011111100: color_data = 12'b111011101110;
20'b00100000110011111101: color_data = 12'b111011101110;
20'b00100000110011111110: color_data = 12'b111011101110;
20'b00100000110011111111: color_data = 12'b111011101110;
20'b00100000110100000000: color_data = 12'b111011101110;
20'b00100000110100000001: color_data = 12'b111011101110;
20'b00100000110100000010: color_data = 12'b111011101110;
20'b00100000110100000100: color_data = 12'b111011101110;
20'b00100000110100000101: color_data = 12'b111011101110;
20'b00100000110100000110: color_data = 12'b111011101110;
20'b00100000110100000111: color_data = 12'b111011101110;
20'b00100000110100001000: color_data = 12'b111011101110;
20'b00100000110100001001: color_data = 12'b111011101110;
20'b00100000110100001010: color_data = 12'b111011101110;
20'b00100000110100001011: color_data = 12'b111011101110;
20'b00100000110100001100: color_data = 12'b111011101110;
20'b00100000110100001101: color_data = 12'b111011101110;
20'b00100000110100100101: color_data = 12'b111011101110;
20'b00100000110100100110: color_data = 12'b111011101110;
20'b00100000110100100111: color_data = 12'b111011101110;
20'b00100000110100101000: color_data = 12'b111011101110;
20'b00100000110100101001: color_data = 12'b111011101110;
20'b00100000110100101010: color_data = 12'b111011101110;
20'b00100000110100101011: color_data = 12'b111011101110;
20'b00100000110100101100: color_data = 12'b111011101110;
20'b00100000110100101101: color_data = 12'b111011101110;
20'b00100000110100101110: color_data = 12'b111011101110;
20'b00100000110101000110: color_data = 12'b111011101110;
20'b00100000110101000111: color_data = 12'b111011101110;
20'b00100000110101001000: color_data = 12'b111011101110;
20'b00100000110101001001: color_data = 12'b111011101110;
20'b00100000110101001010: color_data = 12'b111011101110;
20'b00100000110101001011: color_data = 12'b111011101110;
20'b00100000110101001100: color_data = 12'b111011101110;
20'b00100000110101001101: color_data = 12'b111011101110;
20'b00100000110101001110: color_data = 12'b111011101110;
20'b00100000110101001111: color_data = 12'b111011101110;
20'b00100000110101110010: color_data = 12'b111011101110;
20'b00100000110101110011: color_data = 12'b111011101110;
20'b00100000110101110100: color_data = 12'b111011101110;
20'b00100000110101110101: color_data = 12'b111011101110;
20'b00100000110101110110: color_data = 12'b111011101110;
20'b00100000110101110111: color_data = 12'b111011101110;
20'b00100000110101111000: color_data = 12'b111011101110;
20'b00100000110101111001: color_data = 12'b111011101110;
20'b00100000110101111010: color_data = 12'b111011101110;
20'b00100000110101111011: color_data = 12'b111011101110;
20'b00100000110101111101: color_data = 12'b111011101110;
20'b00100000110101111110: color_data = 12'b111011101110;
20'b00100000110101111111: color_data = 12'b111011101110;
20'b00100000110110000000: color_data = 12'b111011101110;
20'b00100000110110000001: color_data = 12'b111011101110;
20'b00100000110110000010: color_data = 12'b111011101110;
20'b00100000110110000011: color_data = 12'b111011101110;
20'b00100000110110000100: color_data = 12'b111011101110;
20'b00100000110110000101: color_data = 12'b111011101110;
20'b00100000110110000110: color_data = 12'b111011101110;
20'b00100000110110001000: color_data = 12'b111011101110;
20'b00100000110110001001: color_data = 12'b111011101110;
20'b00100000110110001010: color_data = 12'b111011101110;
20'b00100000110110001011: color_data = 12'b111011101110;
20'b00100000110110001100: color_data = 12'b111011101110;
20'b00100000110110001101: color_data = 12'b111011101110;
20'b00100000110110001110: color_data = 12'b111011101110;
20'b00100000110110001111: color_data = 12'b111011101110;
20'b00100000110110010000: color_data = 12'b111011101110;
20'b00100000110110010001: color_data = 12'b111011101110;
20'b00100000110110101001: color_data = 12'b111011101110;
20'b00100000110110101010: color_data = 12'b111011101110;
20'b00100000110110101011: color_data = 12'b111011101110;
20'b00100000110110101100: color_data = 12'b111011101110;
20'b00100000110110101101: color_data = 12'b111011101110;
20'b00100000110110101110: color_data = 12'b111011101110;
20'b00100000110110101111: color_data = 12'b111011101110;
20'b00100000110110110000: color_data = 12'b111011101110;
20'b00100000110110110001: color_data = 12'b111011101110;
20'b00100000110110110010: color_data = 12'b111011101110;
20'b00100001000011001101: color_data = 12'b111011101110;
20'b00100001000011001110: color_data = 12'b111011101110;
20'b00100001000011001111: color_data = 12'b111011101110;
20'b00100001000011010000: color_data = 12'b111011101110;
20'b00100001000011010001: color_data = 12'b111011101110;
20'b00100001000011010010: color_data = 12'b111011101110;
20'b00100001000011010011: color_data = 12'b111011101110;
20'b00100001000011010100: color_data = 12'b111011101110;
20'b00100001000011010101: color_data = 12'b111011101110;
20'b00100001000011010110: color_data = 12'b111011101110;
20'b00100001000011011000: color_data = 12'b111011101110;
20'b00100001000011011001: color_data = 12'b111011101110;
20'b00100001000011011010: color_data = 12'b111011101110;
20'b00100001000011011011: color_data = 12'b111011101110;
20'b00100001000011011100: color_data = 12'b111011101110;
20'b00100001000011011101: color_data = 12'b111011101110;
20'b00100001000011011110: color_data = 12'b111011101110;
20'b00100001000011011111: color_data = 12'b111011101110;
20'b00100001000011100000: color_data = 12'b111011101110;
20'b00100001000011100001: color_data = 12'b111011101110;
20'b00100001000011111001: color_data = 12'b111011101110;
20'b00100001000011111010: color_data = 12'b111011101110;
20'b00100001000011111011: color_data = 12'b111011101110;
20'b00100001000011111100: color_data = 12'b111011101110;
20'b00100001000011111101: color_data = 12'b111011101110;
20'b00100001000011111110: color_data = 12'b111011101110;
20'b00100001000011111111: color_data = 12'b111011101110;
20'b00100001000100000000: color_data = 12'b111011101110;
20'b00100001000100000001: color_data = 12'b111011101110;
20'b00100001000100000010: color_data = 12'b111011101110;
20'b00100001000100000100: color_data = 12'b111011101110;
20'b00100001000100000101: color_data = 12'b111011101110;
20'b00100001000100000110: color_data = 12'b111011101110;
20'b00100001000100000111: color_data = 12'b111011101110;
20'b00100001000100001000: color_data = 12'b111011101110;
20'b00100001000100001001: color_data = 12'b111011101110;
20'b00100001000100001010: color_data = 12'b111011101110;
20'b00100001000100001011: color_data = 12'b111011101110;
20'b00100001000100001100: color_data = 12'b111011101110;
20'b00100001000100001101: color_data = 12'b111011101110;
20'b00100001000100100101: color_data = 12'b111011101110;
20'b00100001000100100110: color_data = 12'b111011101110;
20'b00100001000100100111: color_data = 12'b111011101110;
20'b00100001000100101000: color_data = 12'b111011101110;
20'b00100001000100101001: color_data = 12'b111011101110;
20'b00100001000100101010: color_data = 12'b111011101110;
20'b00100001000100101011: color_data = 12'b111011101110;
20'b00100001000100101100: color_data = 12'b111011101110;
20'b00100001000100101101: color_data = 12'b111011101110;
20'b00100001000100101110: color_data = 12'b111011101110;
20'b00100001000101000110: color_data = 12'b111011101110;
20'b00100001000101000111: color_data = 12'b111011101110;
20'b00100001000101001000: color_data = 12'b111011101110;
20'b00100001000101001001: color_data = 12'b111011101110;
20'b00100001000101001010: color_data = 12'b111011101110;
20'b00100001000101001011: color_data = 12'b111011101110;
20'b00100001000101001100: color_data = 12'b111011101110;
20'b00100001000101001101: color_data = 12'b111011101110;
20'b00100001000101001110: color_data = 12'b111011101110;
20'b00100001000101001111: color_data = 12'b111011101110;
20'b00100001000101110010: color_data = 12'b111011101110;
20'b00100001000101110011: color_data = 12'b111011101110;
20'b00100001000101110100: color_data = 12'b111011101110;
20'b00100001000101110101: color_data = 12'b111011101110;
20'b00100001000101110110: color_data = 12'b111011101110;
20'b00100001000101110111: color_data = 12'b111011101110;
20'b00100001000101111000: color_data = 12'b111011101110;
20'b00100001000101111001: color_data = 12'b111011101110;
20'b00100001000101111010: color_data = 12'b111011101110;
20'b00100001000101111011: color_data = 12'b111011101110;
20'b00100001000101111101: color_data = 12'b111011101110;
20'b00100001000101111110: color_data = 12'b111011101110;
20'b00100001000101111111: color_data = 12'b111011101110;
20'b00100001000110000000: color_data = 12'b111011101110;
20'b00100001000110000001: color_data = 12'b111011101110;
20'b00100001000110000010: color_data = 12'b111011101110;
20'b00100001000110000011: color_data = 12'b111011101110;
20'b00100001000110000100: color_data = 12'b111011101110;
20'b00100001000110000101: color_data = 12'b111011101110;
20'b00100001000110000110: color_data = 12'b111011101110;
20'b00100001000110001000: color_data = 12'b111011101110;
20'b00100001000110001001: color_data = 12'b111011101110;
20'b00100001000110001010: color_data = 12'b111011101110;
20'b00100001000110001011: color_data = 12'b111011101110;
20'b00100001000110001100: color_data = 12'b111011101110;
20'b00100001000110001101: color_data = 12'b111011101110;
20'b00100001000110001110: color_data = 12'b111011101110;
20'b00100001000110001111: color_data = 12'b111011101110;
20'b00100001000110010000: color_data = 12'b111011101110;
20'b00100001000110010001: color_data = 12'b111011101110;
20'b00100001000110101001: color_data = 12'b111011101110;
20'b00100001000110101010: color_data = 12'b111011101110;
20'b00100001000110101011: color_data = 12'b111011101110;
20'b00100001000110101100: color_data = 12'b111011101110;
20'b00100001000110101101: color_data = 12'b111011101110;
20'b00100001000110101110: color_data = 12'b111011101110;
20'b00100001000110101111: color_data = 12'b111011101110;
20'b00100001000110110000: color_data = 12'b111011101110;
20'b00100001000110110001: color_data = 12'b111011101110;
20'b00100001000110110010: color_data = 12'b111011101110;
20'b00100001010011001101: color_data = 12'b111011101110;
20'b00100001010011001110: color_data = 12'b111011101110;
20'b00100001010011001111: color_data = 12'b111011101110;
20'b00100001010011010000: color_data = 12'b111011101110;
20'b00100001010011010001: color_data = 12'b111011101110;
20'b00100001010011010010: color_data = 12'b111011101110;
20'b00100001010011010011: color_data = 12'b111011101110;
20'b00100001010011010100: color_data = 12'b111011101110;
20'b00100001010011010101: color_data = 12'b111011101110;
20'b00100001010011010110: color_data = 12'b111011101110;
20'b00100001010011011000: color_data = 12'b111011101110;
20'b00100001010011011001: color_data = 12'b111011101110;
20'b00100001010011011010: color_data = 12'b111011101110;
20'b00100001010011011011: color_data = 12'b111011101110;
20'b00100001010011011100: color_data = 12'b111011101110;
20'b00100001010011011101: color_data = 12'b111011101110;
20'b00100001010011011110: color_data = 12'b111011101110;
20'b00100001010011011111: color_data = 12'b111011101110;
20'b00100001010011100000: color_data = 12'b111011101110;
20'b00100001010011100001: color_data = 12'b111011101110;
20'b00100001010011111001: color_data = 12'b111011101110;
20'b00100001010011111010: color_data = 12'b111011101110;
20'b00100001010011111011: color_data = 12'b111011101110;
20'b00100001010011111100: color_data = 12'b111011101110;
20'b00100001010011111101: color_data = 12'b111011101110;
20'b00100001010011111110: color_data = 12'b111011101110;
20'b00100001010011111111: color_data = 12'b111011101110;
20'b00100001010100000000: color_data = 12'b111011101110;
20'b00100001010100000001: color_data = 12'b111011101110;
20'b00100001010100000010: color_data = 12'b111011101110;
20'b00100001010100000100: color_data = 12'b111011101110;
20'b00100001010100000101: color_data = 12'b111011101110;
20'b00100001010100000110: color_data = 12'b111011101110;
20'b00100001010100000111: color_data = 12'b111011101110;
20'b00100001010100001000: color_data = 12'b111011101110;
20'b00100001010100001001: color_data = 12'b111011101110;
20'b00100001010100001010: color_data = 12'b111011101110;
20'b00100001010100001011: color_data = 12'b111011101110;
20'b00100001010100001100: color_data = 12'b111011101110;
20'b00100001010100001101: color_data = 12'b111011101110;
20'b00100001010100100101: color_data = 12'b111011101110;
20'b00100001010100100110: color_data = 12'b111011101110;
20'b00100001010100100111: color_data = 12'b111011101110;
20'b00100001010100101000: color_data = 12'b111011101110;
20'b00100001010100101001: color_data = 12'b111011101110;
20'b00100001010100101010: color_data = 12'b111011101110;
20'b00100001010100101011: color_data = 12'b111011101110;
20'b00100001010100101100: color_data = 12'b111011101110;
20'b00100001010100101101: color_data = 12'b111011101110;
20'b00100001010100101110: color_data = 12'b111011101110;
20'b00100001010101000110: color_data = 12'b111011101110;
20'b00100001010101000111: color_data = 12'b111011101110;
20'b00100001010101001000: color_data = 12'b111011101110;
20'b00100001010101001001: color_data = 12'b111011101110;
20'b00100001010101001010: color_data = 12'b111011101110;
20'b00100001010101001011: color_data = 12'b111011101110;
20'b00100001010101001100: color_data = 12'b111011101110;
20'b00100001010101001101: color_data = 12'b111011101110;
20'b00100001010101001110: color_data = 12'b111011101110;
20'b00100001010101001111: color_data = 12'b111011101110;
20'b00100001010101110010: color_data = 12'b111011101110;
20'b00100001010101110011: color_data = 12'b111011101110;
20'b00100001010101110100: color_data = 12'b111011101110;
20'b00100001010101110101: color_data = 12'b111011101110;
20'b00100001010101110110: color_data = 12'b111011101110;
20'b00100001010101110111: color_data = 12'b111011101110;
20'b00100001010101111000: color_data = 12'b111011101110;
20'b00100001010101111001: color_data = 12'b111011101110;
20'b00100001010101111010: color_data = 12'b111011101110;
20'b00100001010101111011: color_data = 12'b111011101110;
20'b00100001010101111101: color_data = 12'b111011101110;
20'b00100001010101111110: color_data = 12'b111011101110;
20'b00100001010101111111: color_data = 12'b111011101110;
20'b00100001010110000000: color_data = 12'b111011101110;
20'b00100001010110000001: color_data = 12'b111011101110;
20'b00100001010110000010: color_data = 12'b111011101110;
20'b00100001010110000011: color_data = 12'b111011101110;
20'b00100001010110000100: color_data = 12'b111011101110;
20'b00100001010110000101: color_data = 12'b111011101110;
20'b00100001010110000110: color_data = 12'b111011101110;
20'b00100001010110001000: color_data = 12'b111011101110;
20'b00100001010110001001: color_data = 12'b111011101110;
20'b00100001010110001010: color_data = 12'b111011101110;
20'b00100001010110001011: color_data = 12'b111011101110;
20'b00100001010110001100: color_data = 12'b111011101110;
20'b00100001010110001101: color_data = 12'b111011101110;
20'b00100001010110001110: color_data = 12'b111011101110;
20'b00100001010110001111: color_data = 12'b111011101110;
20'b00100001010110010000: color_data = 12'b111011101110;
20'b00100001010110010001: color_data = 12'b111011101110;
20'b00100001010110101001: color_data = 12'b111011101110;
20'b00100001010110101010: color_data = 12'b111011101110;
20'b00100001010110101011: color_data = 12'b111011101110;
20'b00100001010110101100: color_data = 12'b111011101110;
20'b00100001010110101101: color_data = 12'b111011101110;
20'b00100001010110101110: color_data = 12'b111011101110;
20'b00100001010110101111: color_data = 12'b111011101110;
20'b00100001010110110000: color_data = 12'b111011101110;
20'b00100001010110110001: color_data = 12'b111011101110;
20'b00100001010110110010: color_data = 12'b111011101110;
20'b00100001100011001101: color_data = 12'b111011101110;
20'b00100001100011001110: color_data = 12'b111011101110;
20'b00100001100011001111: color_data = 12'b111011101110;
20'b00100001100011010000: color_data = 12'b111011101110;
20'b00100001100011010001: color_data = 12'b111011101110;
20'b00100001100011010010: color_data = 12'b111011101110;
20'b00100001100011010011: color_data = 12'b111011101110;
20'b00100001100011010100: color_data = 12'b111011101110;
20'b00100001100011010101: color_data = 12'b111011101110;
20'b00100001100011010110: color_data = 12'b111011101110;
20'b00100001100011011000: color_data = 12'b111011101110;
20'b00100001100011011001: color_data = 12'b111011101110;
20'b00100001100011011010: color_data = 12'b111011101110;
20'b00100001100011011011: color_data = 12'b111011101110;
20'b00100001100011011100: color_data = 12'b111011101110;
20'b00100001100011011101: color_data = 12'b111011101110;
20'b00100001100011011110: color_data = 12'b111011101110;
20'b00100001100011011111: color_data = 12'b111011101110;
20'b00100001100011100000: color_data = 12'b111011101110;
20'b00100001100011100001: color_data = 12'b111011101110;
20'b00100001100011111001: color_data = 12'b111011101110;
20'b00100001100011111010: color_data = 12'b111011101110;
20'b00100001100011111011: color_data = 12'b111011101110;
20'b00100001100011111100: color_data = 12'b111011101110;
20'b00100001100011111101: color_data = 12'b111011101110;
20'b00100001100011111110: color_data = 12'b111011101110;
20'b00100001100011111111: color_data = 12'b111011101110;
20'b00100001100100000000: color_data = 12'b111011101110;
20'b00100001100100000001: color_data = 12'b111011101110;
20'b00100001100100000010: color_data = 12'b111011101110;
20'b00100001100100000100: color_data = 12'b111011101110;
20'b00100001100100000101: color_data = 12'b111011101110;
20'b00100001100100000110: color_data = 12'b111011101110;
20'b00100001100100000111: color_data = 12'b111011101110;
20'b00100001100100001000: color_data = 12'b111011101110;
20'b00100001100100001001: color_data = 12'b111011101110;
20'b00100001100100001010: color_data = 12'b111011101110;
20'b00100001100100001011: color_data = 12'b111011101110;
20'b00100001100100001100: color_data = 12'b111011101110;
20'b00100001100100001101: color_data = 12'b111011101110;
20'b00100001100100100101: color_data = 12'b111011101110;
20'b00100001100100100110: color_data = 12'b111011101110;
20'b00100001100100100111: color_data = 12'b111011101110;
20'b00100001100100101000: color_data = 12'b111011101110;
20'b00100001100100101001: color_data = 12'b111011101110;
20'b00100001100100101010: color_data = 12'b111011101110;
20'b00100001100100101011: color_data = 12'b111011101110;
20'b00100001100100101100: color_data = 12'b111011101110;
20'b00100001100100101101: color_data = 12'b111011101110;
20'b00100001100100101110: color_data = 12'b111011101110;
20'b00100001100101000110: color_data = 12'b111011101110;
20'b00100001100101000111: color_data = 12'b111011101110;
20'b00100001100101001000: color_data = 12'b111011101110;
20'b00100001100101001001: color_data = 12'b111011101110;
20'b00100001100101001010: color_data = 12'b111011101110;
20'b00100001100101001011: color_data = 12'b111011101110;
20'b00100001100101001100: color_data = 12'b111011101110;
20'b00100001100101001101: color_data = 12'b111011101110;
20'b00100001100101001110: color_data = 12'b111011101110;
20'b00100001100101001111: color_data = 12'b111011101110;
20'b00100001100101110010: color_data = 12'b111011101110;
20'b00100001100101110011: color_data = 12'b111011101110;
20'b00100001100101110100: color_data = 12'b111011101110;
20'b00100001100101110101: color_data = 12'b111011101110;
20'b00100001100101110110: color_data = 12'b111011101110;
20'b00100001100101110111: color_data = 12'b111011101110;
20'b00100001100101111000: color_data = 12'b111011101110;
20'b00100001100101111001: color_data = 12'b111011101110;
20'b00100001100101111010: color_data = 12'b111011101110;
20'b00100001100101111011: color_data = 12'b111011101110;
20'b00100001100101111101: color_data = 12'b111011101110;
20'b00100001100101111110: color_data = 12'b111011101110;
20'b00100001100101111111: color_data = 12'b111011101110;
20'b00100001100110000000: color_data = 12'b111011101110;
20'b00100001100110000001: color_data = 12'b111011101110;
20'b00100001100110000010: color_data = 12'b111011101110;
20'b00100001100110000011: color_data = 12'b111011101110;
20'b00100001100110000100: color_data = 12'b111011101110;
20'b00100001100110000101: color_data = 12'b111011101110;
20'b00100001100110000110: color_data = 12'b111011101110;
20'b00100001100110001000: color_data = 12'b111011101110;
20'b00100001100110001001: color_data = 12'b111011101110;
20'b00100001100110001010: color_data = 12'b111011101110;
20'b00100001100110001011: color_data = 12'b111011101110;
20'b00100001100110001100: color_data = 12'b111011101110;
20'b00100001100110001101: color_data = 12'b111011101110;
20'b00100001100110001110: color_data = 12'b111011101110;
20'b00100001100110001111: color_data = 12'b111011101110;
20'b00100001100110010000: color_data = 12'b111011101110;
20'b00100001100110010001: color_data = 12'b111011101110;
20'b00100001100110101001: color_data = 12'b111011101110;
20'b00100001100110101010: color_data = 12'b111011101110;
20'b00100001100110101011: color_data = 12'b111011101110;
20'b00100001100110101100: color_data = 12'b111011101110;
20'b00100001100110101101: color_data = 12'b111011101110;
20'b00100001100110101110: color_data = 12'b111011101110;
20'b00100001100110101111: color_data = 12'b111011101110;
20'b00100001100110110000: color_data = 12'b111011101110;
20'b00100001100110110001: color_data = 12'b111011101110;
20'b00100001100110110010: color_data = 12'b111011101110;
20'b00100001110011001101: color_data = 12'b111011101110;
20'b00100001110011001110: color_data = 12'b111011101110;
20'b00100001110011001111: color_data = 12'b111011101110;
20'b00100001110011010000: color_data = 12'b111011101110;
20'b00100001110011010001: color_data = 12'b111011101110;
20'b00100001110011010010: color_data = 12'b111011101110;
20'b00100001110011010011: color_data = 12'b111011101110;
20'b00100001110011010100: color_data = 12'b111011101110;
20'b00100001110011010101: color_data = 12'b111011101110;
20'b00100001110011010110: color_data = 12'b111011101110;
20'b00100001110011011000: color_data = 12'b111011101110;
20'b00100001110011011001: color_data = 12'b111011101110;
20'b00100001110011011010: color_data = 12'b111011101110;
20'b00100001110011011011: color_data = 12'b111011101110;
20'b00100001110011011100: color_data = 12'b111011101110;
20'b00100001110011011101: color_data = 12'b111011101110;
20'b00100001110011011110: color_data = 12'b111011101110;
20'b00100001110011011111: color_data = 12'b111011101110;
20'b00100001110011100000: color_data = 12'b111011101110;
20'b00100001110011100001: color_data = 12'b111011101110;
20'b00100001110011111001: color_data = 12'b111011101110;
20'b00100001110011111010: color_data = 12'b111011101110;
20'b00100001110011111011: color_data = 12'b111011101110;
20'b00100001110011111100: color_data = 12'b111011101110;
20'b00100001110011111101: color_data = 12'b111011101110;
20'b00100001110011111110: color_data = 12'b111011101110;
20'b00100001110011111111: color_data = 12'b111011101110;
20'b00100001110100000000: color_data = 12'b111011101110;
20'b00100001110100000001: color_data = 12'b111011101110;
20'b00100001110100000010: color_data = 12'b111011101110;
20'b00100001110100000100: color_data = 12'b111011101110;
20'b00100001110100000101: color_data = 12'b111011101110;
20'b00100001110100000110: color_data = 12'b111011101110;
20'b00100001110100000111: color_data = 12'b111011101110;
20'b00100001110100001000: color_data = 12'b111011101110;
20'b00100001110100001001: color_data = 12'b111011101110;
20'b00100001110100001010: color_data = 12'b111011101110;
20'b00100001110100001011: color_data = 12'b111011101110;
20'b00100001110100001100: color_data = 12'b111011101110;
20'b00100001110100001101: color_data = 12'b111011101110;
20'b00100001110100100101: color_data = 12'b111011101110;
20'b00100001110100100110: color_data = 12'b111011101110;
20'b00100001110100100111: color_data = 12'b111011101110;
20'b00100001110100101000: color_data = 12'b111011101110;
20'b00100001110100101001: color_data = 12'b111011101110;
20'b00100001110100101010: color_data = 12'b111011101110;
20'b00100001110100101011: color_data = 12'b111011101110;
20'b00100001110100101100: color_data = 12'b111011101110;
20'b00100001110100101101: color_data = 12'b111011101110;
20'b00100001110100101110: color_data = 12'b111011101110;
20'b00100001110101000110: color_data = 12'b111011101110;
20'b00100001110101000111: color_data = 12'b111011101110;
20'b00100001110101001000: color_data = 12'b111011101110;
20'b00100001110101001001: color_data = 12'b111011101110;
20'b00100001110101001010: color_data = 12'b111011101110;
20'b00100001110101001011: color_data = 12'b111011101110;
20'b00100001110101001100: color_data = 12'b111011101110;
20'b00100001110101001101: color_data = 12'b111011101110;
20'b00100001110101001110: color_data = 12'b111011101110;
20'b00100001110101001111: color_data = 12'b111011101110;
20'b00100001110101110010: color_data = 12'b111011101110;
20'b00100001110101110011: color_data = 12'b111011101110;
20'b00100001110101110100: color_data = 12'b111011101110;
20'b00100001110101110101: color_data = 12'b111011101110;
20'b00100001110101110110: color_data = 12'b111011101110;
20'b00100001110101110111: color_data = 12'b111011101110;
20'b00100001110101111000: color_data = 12'b111011101110;
20'b00100001110101111001: color_data = 12'b111011101110;
20'b00100001110101111010: color_data = 12'b111011101110;
20'b00100001110101111011: color_data = 12'b111011101110;
20'b00100001110101111101: color_data = 12'b111011101110;
20'b00100001110101111110: color_data = 12'b111011101110;
20'b00100001110101111111: color_data = 12'b111011101110;
20'b00100001110110000000: color_data = 12'b111011101110;
20'b00100001110110000001: color_data = 12'b111011101110;
20'b00100001110110000010: color_data = 12'b111011101110;
20'b00100001110110000011: color_data = 12'b111011101110;
20'b00100001110110000100: color_data = 12'b111011101110;
20'b00100001110110000101: color_data = 12'b111011101110;
20'b00100001110110000110: color_data = 12'b111011101110;
20'b00100001110110001000: color_data = 12'b111011101110;
20'b00100001110110001001: color_data = 12'b111011101110;
20'b00100001110110001010: color_data = 12'b111011101110;
20'b00100001110110001011: color_data = 12'b111011101110;
20'b00100001110110001100: color_data = 12'b111011101110;
20'b00100001110110001101: color_data = 12'b111011101110;
20'b00100001110110001110: color_data = 12'b111011101110;
20'b00100001110110001111: color_data = 12'b111011101110;
20'b00100001110110010000: color_data = 12'b111011101110;
20'b00100001110110010001: color_data = 12'b111011101110;
20'b00100001110110101001: color_data = 12'b111011101110;
20'b00100001110110101010: color_data = 12'b111011101110;
20'b00100001110110101011: color_data = 12'b111011101110;
20'b00100001110110101100: color_data = 12'b111011101110;
20'b00100001110110101101: color_data = 12'b111011101110;
20'b00100001110110101110: color_data = 12'b111011101110;
20'b00100001110110101111: color_data = 12'b111011101110;
20'b00100001110110110000: color_data = 12'b111011101110;
20'b00100001110110110001: color_data = 12'b111011101110;
20'b00100001110110110010: color_data = 12'b111011101110;
20'b00100010010010010110: color_data = 12'b111011101110;
20'b00100010010010010111: color_data = 12'b111011101110;
20'b00100010010010011000: color_data = 12'b111011101110;
20'b00100010010010011001: color_data = 12'b111011101110;
20'b00100010010010011010: color_data = 12'b111011101110;
20'b00100010010010011011: color_data = 12'b111011101110;
20'b00100010010010011100: color_data = 12'b111011101110;
20'b00100010010010011101: color_data = 12'b111011101110;
20'b00100010010010011110: color_data = 12'b111011101110;
20'b00100010010010011111: color_data = 12'b111011101110;
20'b00100010010010100001: color_data = 12'b111011101110;
20'b00100010010010100010: color_data = 12'b111011101110;
20'b00100010010010100011: color_data = 12'b111011101110;
20'b00100010010010100100: color_data = 12'b111011101110;
20'b00100010010010100101: color_data = 12'b111011101110;
20'b00100010010010100110: color_data = 12'b111011101110;
20'b00100010010010100111: color_data = 12'b111011101110;
20'b00100010010010101000: color_data = 12'b111011101110;
20'b00100010010010101001: color_data = 12'b111011101110;
20'b00100010010010101010: color_data = 12'b111011101110;
20'b00100010010011101110: color_data = 12'b111011101110;
20'b00100010010011101111: color_data = 12'b111011101110;
20'b00100010010011110000: color_data = 12'b111011101110;
20'b00100010010011110001: color_data = 12'b111011101110;
20'b00100010010011110010: color_data = 12'b111011101110;
20'b00100010010011110011: color_data = 12'b111011101110;
20'b00100010010011110100: color_data = 12'b111011101110;
20'b00100010010011110101: color_data = 12'b111011101110;
20'b00100010010011110110: color_data = 12'b111011101110;
20'b00100010010011110111: color_data = 12'b111011101110;
20'b00100010010011111001: color_data = 12'b111011101110;
20'b00100010010011111010: color_data = 12'b111011101110;
20'b00100010010011111011: color_data = 12'b111011101110;
20'b00100010010011111100: color_data = 12'b111011101110;
20'b00100010010011111101: color_data = 12'b111011101110;
20'b00100010010011111110: color_data = 12'b111011101110;
20'b00100010010011111111: color_data = 12'b111011101110;
20'b00100010010100000000: color_data = 12'b111011101110;
20'b00100010010100000001: color_data = 12'b111011101110;
20'b00100010010100000010: color_data = 12'b111011101110;
20'b00100010010100100101: color_data = 12'b111011101110;
20'b00100010010100100110: color_data = 12'b111011101110;
20'b00100010010100100111: color_data = 12'b111011101110;
20'b00100010010100101000: color_data = 12'b111011101110;
20'b00100010010100101001: color_data = 12'b111011101110;
20'b00100010010100101010: color_data = 12'b111011101110;
20'b00100010010100101011: color_data = 12'b111011101110;
20'b00100010010100101100: color_data = 12'b111011101110;
20'b00100010010100101101: color_data = 12'b111011101110;
20'b00100010010100101110: color_data = 12'b111011101110;
20'b00100010010100110000: color_data = 12'b111011101110;
20'b00100010010100110001: color_data = 12'b111011101110;
20'b00100010010100110010: color_data = 12'b111011101110;
20'b00100010010100110011: color_data = 12'b111011101110;
20'b00100010010100110100: color_data = 12'b111011101110;
20'b00100010010100110101: color_data = 12'b111011101110;
20'b00100010010100110110: color_data = 12'b111011101110;
20'b00100010010100110111: color_data = 12'b111011101110;
20'b00100010010100111000: color_data = 12'b111011101110;
20'b00100010010100111001: color_data = 12'b111011101110;
20'b00100010010101000110: color_data = 12'b111011101110;
20'b00100010010101000111: color_data = 12'b111011101110;
20'b00100010010101001000: color_data = 12'b111011101110;
20'b00100010010101001001: color_data = 12'b111011101110;
20'b00100010010101001010: color_data = 12'b111011101110;
20'b00100010010101001011: color_data = 12'b111011101110;
20'b00100010010101001100: color_data = 12'b111011101110;
20'b00100010010101001101: color_data = 12'b111011101110;
20'b00100010010101001110: color_data = 12'b111011101110;
20'b00100010010101001111: color_data = 12'b111011101110;
20'b00100010010101010001: color_data = 12'b111011101110;
20'b00100010010101010010: color_data = 12'b111011101110;
20'b00100010010101010011: color_data = 12'b111011101110;
20'b00100010010101010100: color_data = 12'b111011101110;
20'b00100010010101010101: color_data = 12'b111011101110;
20'b00100010010101010110: color_data = 12'b111011101110;
20'b00100010010101010111: color_data = 12'b111011101110;
20'b00100010010101011000: color_data = 12'b111011101110;
20'b00100010010101011001: color_data = 12'b111011101110;
20'b00100010010101011010: color_data = 12'b111011101110;
20'b00100010010101011100: color_data = 12'b111011101110;
20'b00100010010101011101: color_data = 12'b111011101110;
20'b00100010010101011110: color_data = 12'b111011101110;
20'b00100010010101011111: color_data = 12'b111011101110;
20'b00100010010101100000: color_data = 12'b111011101110;
20'b00100010010101100001: color_data = 12'b111011101110;
20'b00100010010101100010: color_data = 12'b111011101110;
20'b00100010010101100011: color_data = 12'b111011101110;
20'b00100010010101100100: color_data = 12'b111011101110;
20'b00100010010101100101: color_data = 12'b111011101110;
20'b00100010010101100111: color_data = 12'b111011101110;
20'b00100010010101101000: color_data = 12'b111011101110;
20'b00100010010101101001: color_data = 12'b111011101110;
20'b00100010010101101010: color_data = 12'b111011101110;
20'b00100010010101101011: color_data = 12'b111011101110;
20'b00100010010101101100: color_data = 12'b111011101110;
20'b00100010010101101101: color_data = 12'b111011101110;
20'b00100010010101101110: color_data = 12'b111011101110;
20'b00100010010101101111: color_data = 12'b111011101110;
20'b00100010010101110000: color_data = 12'b111011101110;
20'b00100010010101110010: color_data = 12'b111011101110;
20'b00100010010101110011: color_data = 12'b111011101110;
20'b00100010010101110100: color_data = 12'b111011101110;
20'b00100010010101110101: color_data = 12'b111011101110;
20'b00100010010101110110: color_data = 12'b111011101110;
20'b00100010010101110111: color_data = 12'b111011101110;
20'b00100010010101111000: color_data = 12'b111011101110;
20'b00100010010101111001: color_data = 12'b111011101110;
20'b00100010010101111010: color_data = 12'b111011101110;
20'b00100010010101111011: color_data = 12'b111011101110;
20'b00100010010101111101: color_data = 12'b111011101110;
20'b00100010010101111110: color_data = 12'b111011101110;
20'b00100010010101111111: color_data = 12'b111011101110;
20'b00100010010110000000: color_data = 12'b111011101110;
20'b00100010010110000001: color_data = 12'b111011101110;
20'b00100010010110000010: color_data = 12'b111011101110;
20'b00100010010110000011: color_data = 12'b111011101110;
20'b00100010010110000100: color_data = 12'b111011101110;
20'b00100010010110000101: color_data = 12'b111011101110;
20'b00100010010110000110: color_data = 12'b111011101110;
20'b00100010010110001000: color_data = 12'b111011101110;
20'b00100010010110001001: color_data = 12'b111011101110;
20'b00100010010110001010: color_data = 12'b111011101110;
20'b00100010010110001011: color_data = 12'b111011101110;
20'b00100010010110001100: color_data = 12'b111011101110;
20'b00100010010110001101: color_data = 12'b111011101110;
20'b00100010010110001110: color_data = 12'b111011101110;
20'b00100010010110001111: color_data = 12'b111011101110;
20'b00100010010110010000: color_data = 12'b111011101110;
20'b00100010010110010001: color_data = 12'b111011101110;
20'b00100010010110101001: color_data = 12'b111011101110;
20'b00100010010110101010: color_data = 12'b111011101110;
20'b00100010010110101011: color_data = 12'b111011101110;
20'b00100010010110101100: color_data = 12'b111011101110;
20'b00100010010110101101: color_data = 12'b111011101110;
20'b00100010010110101110: color_data = 12'b111011101110;
20'b00100010010110101111: color_data = 12'b111011101110;
20'b00100010010110110000: color_data = 12'b111011101110;
20'b00100010010110110001: color_data = 12'b111011101110;
20'b00100010010110110010: color_data = 12'b111011101110;
20'b00100010100010010110: color_data = 12'b111011101110;
20'b00100010100010010111: color_data = 12'b111011101110;
20'b00100010100010011000: color_data = 12'b111011101110;
20'b00100010100010011001: color_data = 12'b111011101110;
20'b00100010100010011010: color_data = 12'b111011101110;
20'b00100010100010011011: color_data = 12'b111011101110;
20'b00100010100010011100: color_data = 12'b111011101110;
20'b00100010100010011101: color_data = 12'b111011101110;
20'b00100010100010011110: color_data = 12'b111011101110;
20'b00100010100010011111: color_data = 12'b111011101110;
20'b00100010100010100001: color_data = 12'b111011101110;
20'b00100010100010100010: color_data = 12'b111011101110;
20'b00100010100010100011: color_data = 12'b111011101110;
20'b00100010100010100100: color_data = 12'b111011101110;
20'b00100010100010100101: color_data = 12'b111011101110;
20'b00100010100010100110: color_data = 12'b111011101110;
20'b00100010100010100111: color_data = 12'b111011101110;
20'b00100010100010101000: color_data = 12'b111011101110;
20'b00100010100010101001: color_data = 12'b111011101110;
20'b00100010100010101010: color_data = 12'b111011101110;
20'b00100010100011101110: color_data = 12'b111011101110;
20'b00100010100011101111: color_data = 12'b111011101110;
20'b00100010100011110000: color_data = 12'b111011101110;
20'b00100010100011110001: color_data = 12'b111011101110;
20'b00100010100011110010: color_data = 12'b111011101110;
20'b00100010100011110011: color_data = 12'b111011101110;
20'b00100010100011110100: color_data = 12'b111011101110;
20'b00100010100011110101: color_data = 12'b111011101110;
20'b00100010100011110110: color_data = 12'b111011101110;
20'b00100010100011110111: color_data = 12'b111011101110;
20'b00100010100011111001: color_data = 12'b111011101110;
20'b00100010100011111010: color_data = 12'b111011101110;
20'b00100010100011111011: color_data = 12'b111011101110;
20'b00100010100011111100: color_data = 12'b111011101110;
20'b00100010100011111101: color_data = 12'b111011101110;
20'b00100010100011111110: color_data = 12'b111011101110;
20'b00100010100011111111: color_data = 12'b111011101110;
20'b00100010100100000000: color_data = 12'b111011101110;
20'b00100010100100000001: color_data = 12'b111011101110;
20'b00100010100100000010: color_data = 12'b111011101110;
20'b00100010100100100101: color_data = 12'b111011101110;
20'b00100010100100100110: color_data = 12'b111011101110;
20'b00100010100100100111: color_data = 12'b111011101110;
20'b00100010100100101000: color_data = 12'b111011101110;
20'b00100010100100101001: color_data = 12'b111011101110;
20'b00100010100100101010: color_data = 12'b111011101110;
20'b00100010100100101011: color_data = 12'b111011101110;
20'b00100010100100101100: color_data = 12'b111011101110;
20'b00100010100100101101: color_data = 12'b111011101110;
20'b00100010100100101110: color_data = 12'b111011101110;
20'b00100010100100110000: color_data = 12'b111011101110;
20'b00100010100100110001: color_data = 12'b111011101110;
20'b00100010100100110010: color_data = 12'b111011101110;
20'b00100010100100110011: color_data = 12'b111011101110;
20'b00100010100100110100: color_data = 12'b111011101110;
20'b00100010100100110101: color_data = 12'b111011101110;
20'b00100010100100110110: color_data = 12'b111011101110;
20'b00100010100100110111: color_data = 12'b111011101110;
20'b00100010100100111000: color_data = 12'b111011101110;
20'b00100010100100111001: color_data = 12'b111011101110;
20'b00100010100101000110: color_data = 12'b111011101110;
20'b00100010100101000111: color_data = 12'b111011101110;
20'b00100010100101001000: color_data = 12'b111011101110;
20'b00100010100101001001: color_data = 12'b111011101110;
20'b00100010100101001010: color_data = 12'b111011101110;
20'b00100010100101001011: color_data = 12'b111011101110;
20'b00100010100101001100: color_data = 12'b111011101110;
20'b00100010100101001101: color_data = 12'b111011101110;
20'b00100010100101001110: color_data = 12'b111011101110;
20'b00100010100101001111: color_data = 12'b111011101110;
20'b00100010100101010001: color_data = 12'b111011101110;
20'b00100010100101010010: color_data = 12'b111011101110;
20'b00100010100101010011: color_data = 12'b111011101110;
20'b00100010100101010100: color_data = 12'b111011101110;
20'b00100010100101010101: color_data = 12'b111011101110;
20'b00100010100101010110: color_data = 12'b111011101110;
20'b00100010100101010111: color_data = 12'b111011101110;
20'b00100010100101011000: color_data = 12'b111011101110;
20'b00100010100101011001: color_data = 12'b111011101110;
20'b00100010100101011010: color_data = 12'b111011101110;
20'b00100010100101011100: color_data = 12'b111011101110;
20'b00100010100101011101: color_data = 12'b111011101110;
20'b00100010100101011110: color_data = 12'b111011101110;
20'b00100010100101011111: color_data = 12'b111011101110;
20'b00100010100101100000: color_data = 12'b111011101110;
20'b00100010100101100001: color_data = 12'b111011101110;
20'b00100010100101100010: color_data = 12'b111011101110;
20'b00100010100101100011: color_data = 12'b111011101110;
20'b00100010100101100100: color_data = 12'b111011101110;
20'b00100010100101100101: color_data = 12'b111011101110;
20'b00100010100101100111: color_data = 12'b111011101110;
20'b00100010100101101000: color_data = 12'b111011101110;
20'b00100010100101101001: color_data = 12'b111011101110;
20'b00100010100101101010: color_data = 12'b111011101110;
20'b00100010100101101011: color_data = 12'b111011101110;
20'b00100010100101101100: color_data = 12'b111011101110;
20'b00100010100101101101: color_data = 12'b111011101110;
20'b00100010100101101110: color_data = 12'b111011101110;
20'b00100010100101101111: color_data = 12'b111011101110;
20'b00100010100101110000: color_data = 12'b111011101110;
20'b00100010100101110010: color_data = 12'b111011101110;
20'b00100010100101110011: color_data = 12'b111011101110;
20'b00100010100101110100: color_data = 12'b111011101110;
20'b00100010100101110101: color_data = 12'b111011101110;
20'b00100010100101110110: color_data = 12'b111011101110;
20'b00100010100101110111: color_data = 12'b111011101110;
20'b00100010100101111000: color_data = 12'b111011101110;
20'b00100010100101111001: color_data = 12'b111011101110;
20'b00100010100101111010: color_data = 12'b111011101110;
20'b00100010100101111011: color_data = 12'b111011101110;
20'b00100010100101111101: color_data = 12'b111011101110;
20'b00100010100101111110: color_data = 12'b111011101110;
20'b00100010100101111111: color_data = 12'b111011101110;
20'b00100010100110000000: color_data = 12'b111011101110;
20'b00100010100110000001: color_data = 12'b111011101110;
20'b00100010100110000010: color_data = 12'b111011101110;
20'b00100010100110000011: color_data = 12'b111011101110;
20'b00100010100110000100: color_data = 12'b111011101110;
20'b00100010100110000101: color_data = 12'b111011101110;
20'b00100010100110000110: color_data = 12'b111011101110;
20'b00100010100110001000: color_data = 12'b111011101110;
20'b00100010100110001001: color_data = 12'b111011101110;
20'b00100010100110001010: color_data = 12'b111011101110;
20'b00100010100110001011: color_data = 12'b111011101110;
20'b00100010100110001100: color_data = 12'b111011101110;
20'b00100010100110001101: color_data = 12'b111011101110;
20'b00100010100110001110: color_data = 12'b111011101110;
20'b00100010100110001111: color_data = 12'b111011101110;
20'b00100010100110010000: color_data = 12'b111011101110;
20'b00100010100110010001: color_data = 12'b111011101110;
20'b00100010100110101001: color_data = 12'b111011101110;
20'b00100010100110101010: color_data = 12'b111011101110;
20'b00100010100110101011: color_data = 12'b111011101110;
20'b00100010100110101100: color_data = 12'b111011101110;
20'b00100010100110101101: color_data = 12'b111011101110;
20'b00100010100110101110: color_data = 12'b111011101110;
20'b00100010100110101111: color_data = 12'b111011101110;
20'b00100010100110110000: color_data = 12'b111011101110;
20'b00100010100110110001: color_data = 12'b111011101110;
20'b00100010100110110010: color_data = 12'b111011101110;
20'b00100010110010010110: color_data = 12'b111011101110;
20'b00100010110010010111: color_data = 12'b111011101110;
20'b00100010110010011000: color_data = 12'b111011101110;
20'b00100010110010011001: color_data = 12'b111011101110;
20'b00100010110010011010: color_data = 12'b111011101110;
20'b00100010110010011011: color_data = 12'b111011101110;
20'b00100010110010011100: color_data = 12'b111011101110;
20'b00100010110010011101: color_data = 12'b111011101110;
20'b00100010110010011110: color_data = 12'b111011101110;
20'b00100010110010011111: color_data = 12'b111011101110;
20'b00100010110010100001: color_data = 12'b111011101110;
20'b00100010110010100010: color_data = 12'b111011101110;
20'b00100010110010100011: color_data = 12'b111011101110;
20'b00100010110010100100: color_data = 12'b111011101110;
20'b00100010110010100101: color_data = 12'b111011101110;
20'b00100010110010100110: color_data = 12'b111011101110;
20'b00100010110010100111: color_data = 12'b111011101110;
20'b00100010110010101000: color_data = 12'b111011101110;
20'b00100010110010101001: color_data = 12'b111011101110;
20'b00100010110010101010: color_data = 12'b111011101110;
20'b00100010110011101110: color_data = 12'b111011101110;
20'b00100010110011101111: color_data = 12'b111011101110;
20'b00100010110011110000: color_data = 12'b111011101110;
20'b00100010110011110001: color_data = 12'b111011101110;
20'b00100010110011110010: color_data = 12'b111011101110;
20'b00100010110011110011: color_data = 12'b111011101110;
20'b00100010110011110100: color_data = 12'b111011101110;
20'b00100010110011110101: color_data = 12'b111011101110;
20'b00100010110011110110: color_data = 12'b111011101110;
20'b00100010110011110111: color_data = 12'b111011101110;
20'b00100010110011111001: color_data = 12'b111011101110;
20'b00100010110011111010: color_data = 12'b111011101110;
20'b00100010110011111011: color_data = 12'b111011101110;
20'b00100010110011111100: color_data = 12'b111011101110;
20'b00100010110011111101: color_data = 12'b111011101110;
20'b00100010110011111110: color_data = 12'b111011101110;
20'b00100010110011111111: color_data = 12'b111011101110;
20'b00100010110100000000: color_data = 12'b111011101110;
20'b00100010110100000001: color_data = 12'b111011101110;
20'b00100010110100000010: color_data = 12'b111011101110;
20'b00100010110100100101: color_data = 12'b111011101110;
20'b00100010110100100110: color_data = 12'b111011101110;
20'b00100010110100100111: color_data = 12'b111011101110;
20'b00100010110100101000: color_data = 12'b111011101110;
20'b00100010110100101001: color_data = 12'b111011101110;
20'b00100010110100101010: color_data = 12'b111011101110;
20'b00100010110100101011: color_data = 12'b111011101110;
20'b00100010110100101100: color_data = 12'b111011101110;
20'b00100010110100101101: color_data = 12'b111011101110;
20'b00100010110100101110: color_data = 12'b111011101110;
20'b00100010110100110000: color_data = 12'b111011101110;
20'b00100010110100110001: color_data = 12'b111011101110;
20'b00100010110100110010: color_data = 12'b111011101110;
20'b00100010110100110011: color_data = 12'b111011101110;
20'b00100010110100110100: color_data = 12'b111011101110;
20'b00100010110100110101: color_data = 12'b111011101110;
20'b00100010110100110110: color_data = 12'b111011101110;
20'b00100010110100110111: color_data = 12'b111011101110;
20'b00100010110100111000: color_data = 12'b111011101110;
20'b00100010110100111001: color_data = 12'b111011101110;
20'b00100010110101000110: color_data = 12'b111011101110;
20'b00100010110101000111: color_data = 12'b111011101110;
20'b00100010110101001000: color_data = 12'b111011101110;
20'b00100010110101001001: color_data = 12'b111011101110;
20'b00100010110101001010: color_data = 12'b111011101110;
20'b00100010110101001011: color_data = 12'b111011101110;
20'b00100010110101001100: color_data = 12'b111011101110;
20'b00100010110101001101: color_data = 12'b111011101110;
20'b00100010110101001110: color_data = 12'b111011101110;
20'b00100010110101001111: color_data = 12'b111011101110;
20'b00100010110101010001: color_data = 12'b111011101110;
20'b00100010110101010010: color_data = 12'b111011101110;
20'b00100010110101010011: color_data = 12'b111011101110;
20'b00100010110101010100: color_data = 12'b111011101110;
20'b00100010110101010101: color_data = 12'b111011101110;
20'b00100010110101010110: color_data = 12'b111011101110;
20'b00100010110101010111: color_data = 12'b111011101110;
20'b00100010110101011000: color_data = 12'b111011101110;
20'b00100010110101011001: color_data = 12'b111011101110;
20'b00100010110101011010: color_data = 12'b111011101110;
20'b00100010110101011100: color_data = 12'b111011101110;
20'b00100010110101011101: color_data = 12'b111011101110;
20'b00100010110101011110: color_data = 12'b111011101110;
20'b00100010110101011111: color_data = 12'b111011101110;
20'b00100010110101100000: color_data = 12'b111011101110;
20'b00100010110101100001: color_data = 12'b111011101110;
20'b00100010110101100010: color_data = 12'b111011101110;
20'b00100010110101100011: color_data = 12'b111011101110;
20'b00100010110101100100: color_data = 12'b111011101110;
20'b00100010110101100101: color_data = 12'b111011101110;
20'b00100010110101100111: color_data = 12'b111011101110;
20'b00100010110101101000: color_data = 12'b111011101110;
20'b00100010110101101001: color_data = 12'b111011101110;
20'b00100010110101101010: color_data = 12'b111011101110;
20'b00100010110101101011: color_data = 12'b111011101110;
20'b00100010110101101100: color_data = 12'b111011101110;
20'b00100010110101101101: color_data = 12'b111011101110;
20'b00100010110101101110: color_data = 12'b111011101110;
20'b00100010110101101111: color_data = 12'b111011101110;
20'b00100010110101110000: color_data = 12'b111011101110;
20'b00100010110101110010: color_data = 12'b111011101110;
20'b00100010110101110011: color_data = 12'b111011101110;
20'b00100010110101110100: color_data = 12'b111011101110;
20'b00100010110101110101: color_data = 12'b111011101110;
20'b00100010110101110110: color_data = 12'b111011101110;
20'b00100010110101110111: color_data = 12'b111011101110;
20'b00100010110101111000: color_data = 12'b111011101110;
20'b00100010110101111001: color_data = 12'b111011101110;
20'b00100010110101111010: color_data = 12'b111011101110;
20'b00100010110101111011: color_data = 12'b111011101110;
20'b00100010110101111101: color_data = 12'b111011101110;
20'b00100010110101111110: color_data = 12'b111011101110;
20'b00100010110101111111: color_data = 12'b111011101110;
20'b00100010110110000000: color_data = 12'b111011101110;
20'b00100010110110000001: color_data = 12'b111011101110;
20'b00100010110110000010: color_data = 12'b111011101110;
20'b00100010110110000011: color_data = 12'b111011101110;
20'b00100010110110000100: color_data = 12'b111011101110;
20'b00100010110110000101: color_data = 12'b111011101110;
20'b00100010110110000110: color_data = 12'b111011101110;
20'b00100010110110001000: color_data = 12'b111011101110;
20'b00100010110110001001: color_data = 12'b111011101110;
20'b00100010110110001010: color_data = 12'b111011101110;
20'b00100010110110001011: color_data = 12'b111011101110;
20'b00100010110110001100: color_data = 12'b111011101110;
20'b00100010110110001101: color_data = 12'b111011101110;
20'b00100010110110001110: color_data = 12'b111011101110;
20'b00100010110110001111: color_data = 12'b111011101110;
20'b00100010110110010000: color_data = 12'b111011101110;
20'b00100010110110010001: color_data = 12'b111011101110;
20'b00100010110110101001: color_data = 12'b111011101110;
20'b00100010110110101010: color_data = 12'b111011101110;
20'b00100010110110101011: color_data = 12'b111011101110;
20'b00100010110110101100: color_data = 12'b111011101110;
20'b00100010110110101101: color_data = 12'b111011101110;
20'b00100010110110101110: color_data = 12'b111011101110;
20'b00100010110110101111: color_data = 12'b111011101110;
20'b00100010110110110000: color_data = 12'b111011101110;
20'b00100010110110110001: color_data = 12'b111011101110;
20'b00100010110110110010: color_data = 12'b111011101110;
20'b00100011000010010110: color_data = 12'b111011101110;
20'b00100011000010010111: color_data = 12'b111011101110;
20'b00100011000010011000: color_data = 12'b111011101110;
20'b00100011000010011001: color_data = 12'b111011101110;
20'b00100011000010011010: color_data = 12'b111011101110;
20'b00100011000010011011: color_data = 12'b111011101110;
20'b00100011000010011100: color_data = 12'b111011101110;
20'b00100011000010011101: color_data = 12'b111011101110;
20'b00100011000010011110: color_data = 12'b111011101110;
20'b00100011000010011111: color_data = 12'b111011101110;
20'b00100011000010100001: color_data = 12'b111011101110;
20'b00100011000010100010: color_data = 12'b111011101110;
20'b00100011000010100011: color_data = 12'b111011101110;
20'b00100011000010100100: color_data = 12'b111011101110;
20'b00100011000010100101: color_data = 12'b111011101110;
20'b00100011000010100110: color_data = 12'b111011101110;
20'b00100011000010100111: color_data = 12'b111011101110;
20'b00100011000010101000: color_data = 12'b111011101110;
20'b00100011000010101001: color_data = 12'b111011101110;
20'b00100011000010101010: color_data = 12'b111011101110;
20'b00100011000011101110: color_data = 12'b111011101110;
20'b00100011000011101111: color_data = 12'b111011101110;
20'b00100011000011110000: color_data = 12'b111011101110;
20'b00100011000011110001: color_data = 12'b111011101110;
20'b00100011000011110010: color_data = 12'b111011101110;
20'b00100011000011110011: color_data = 12'b111011101110;
20'b00100011000011110100: color_data = 12'b111011101110;
20'b00100011000011110101: color_data = 12'b111011101110;
20'b00100011000011110110: color_data = 12'b111011101110;
20'b00100011000011110111: color_data = 12'b111011101110;
20'b00100011000011111001: color_data = 12'b111011101110;
20'b00100011000011111010: color_data = 12'b111011101110;
20'b00100011000011111011: color_data = 12'b111011101110;
20'b00100011000011111100: color_data = 12'b111011101110;
20'b00100011000011111101: color_data = 12'b111011101110;
20'b00100011000011111110: color_data = 12'b111011101110;
20'b00100011000011111111: color_data = 12'b111011101110;
20'b00100011000100000000: color_data = 12'b111011101110;
20'b00100011000100000001: color_data = 12'b111011101110;
20'b00100011000100000010: color_data = 12'b111011101110;
20'b00100011000100100101: color_data = 12'b111011101110;
20'b00100011000100100110: color_data = 12'b111011101110;
20'b00100011000100100111: color_data = 12'b111011101110;
20'b00100011000100101000: color_data = 12'b111011101110;
20'b00100011000100101001: color_data = 12'b111011101110;
20'b00100011000100101010: color_data = 12'b111011101110;
20'b00100011000100101011: color_data = 12'b111011101110;
20'b00100011000100101100: color_data = 12'b111011101110;
20'b00100011000100101101: color_data = 12'b111011101110;
20'b00100011000100101110: color_data = 12'b111011101110;
20'b00100011000100110000: color_data = 12'b111011101110;
20'b00100011000100110001: color_data = 12'b111011101110;
20'b00100011000100110010: color_data = 12'b111011101110;
20'b00100011000100110011: color_data = 12'b111011101110;
20'b00100011000100110100: color_data = 12'b111011101110;
20'b00100011000100110101: color_data = 12'b111011101110;
20'b00100011000100110110: color_data = 12'b111011101110;
20'b00100011000100110111: color_data = 12'b111011101110;
20'b00100011000100111000: color_data = 12'b111011101110;
20'b00100011000100111001: color_data = 12'b111011101110;
20'b00100011000101000110: color_data = 12'b111011101110;
20'b00100011000101000111: color_data = 12'b111011101110;
20'b00100011000101001000: color_data = 12'b111011101110;
20'b00100011000101001001: color_data = 12'b111011101110;
20'b00100011000101001010: color_data = 12'b111011101110;
20'b00100011000101001011: color_data = 12'b111011101110;
20'b00100011000101001100: color_data = 12'b111011101110;
20'b00100011000101001101: color_data = 12'b111011101110;
20'b00100011000101001110: color_data = 12'b111011101110;
20'b00100011000101001111: color_data = 12'b111011101110;
20'b00100011000101010001: color_data = 12'b111011101110;
20'b00100011000101010010: color_data = 12'b111011101110;
20'b00100011000101010011: color_data = 12'b111011101110;
20'b00100011000101010100: color_data = 12'b111011101110;
20'b00100011000101010101: color_data = 12'b111011101110;
20'b00100011000101010110: color_data = 12'b111011101110;
20'b00100011000101010111: color_data = 12'b111011101110;
20'b00100011000101011000: color_data = 12'b111011101110;
20'b00100011000101011001: color_data = 12'b111011101110;
20'b00100011000101011010: color_data = 12'b111011101110;
20'b00100011000101011100: color_data = 12'b111011101110;
20'b00100011000101011101: color_data = 12'b111011101110;
20'b00100011000101011110: color_data = 12'b111011101110;
20'b00100011000101011111: color_data = 12'b111011101110;
20'b00100011000101100000: color_data = 12'b111011101110;
20'b00100011000101100001: color_data = 12'b111011101110;
20'b00100011000101100010: color_data = 12'b111011101110;
20'b00100011000101100011: color_data = 12'b111011101110;
20'b00100011000101100100: color_data = 12'b111011101110;
20'b00100011000101100101: color_data = 12'b111011101110;
20'b00100011000101100111: color_data = 12'b111011101110;
20'b00100011000101101000: color_data = 12'b111011101110;
20'b00100011000101101001: color_data = 12'b111011101110;
20'b00100011000101101010: color_data = 12'b111011101110;
20'b00100011000101101011: color_data = 12'b111011101110;
20'b00100011000101101100: color_data = 12'b111011101110;
20'b00100011000101101101: color_data = 12'b111011101110;
20'b00100011000101101110: color_data = 12'b111011101110;
20'b00100011000101101111: color_data = 12'b111011101110;
20'b00100011000101110000: color_data = 12'b111011101110;
20'b00100011000101110010: color_data = 12'b111011101110;
20'b00100011000101110011: color_data = 12'b111011101110;
20'b00100011000101110100: color_data = 12'b111011101110;
20'b00100011000101110101: color_data = 12'b111011101110;
20'b00100011000101110110: color_data = 12'b111011101110;
20'b00100011000101110111: color_data = 12'b111011101110;
20'b00100011000101111000: color_data = 12'b111011101110;
20'b00100011000101111001: color_data = 12'b111011101110;
20'b00100011000101111010: color_data = 12'b111011101110;
20'b00100011000101111011: color_data = 12'b111011101110;
20'b00100011000101111101: color_data = 12'b111011101110;
20'b00100011000101111110: color_data = 12'b111011101110;
20'b00100011000101111111: color_data = 12'b111011101110;
20'b00100011000110000000: color_data = 12'b111011101110;
20'b00100011000110000001: color_data = 12'b111011101110;
20'b00100011000110000010: color_data = 12'b111011101110;
20'b00100011000110000011: color_data = 12'b111011101110;
20'b00100011000110000100: color_data = 12'b111011101110;
20'b00100011000110000101: color_data = 12'b111011101110;
20'b00100011000110000110: color_data = 12'b111011101110;
20'b00100011000110001000: color_data = 12'b111011101110;
20'b00100011000110001001: color_data = 12'b111011101110;
20'b00100011000110001010: color_data = 12'b111011101110;
20'b00100011000110001011: color_data = 12'b111011101110;
20'b00100011000110001100: color_data = 12'b111011101110;
20'b00100011000110001101: color_data = 12'b111011101110;
20'b00100011000110001110: color_data = 12'b111011101110;
20'b00100011000110001111: color_data = 12'b111011101110;
20'b00100011000110010000: color_data = 12'b111011101110;
20'b00100011000110010001: color_data = 12'b111011101110;
20'b00100011000110101001: color_data = 12'b111011101110;
20'b00100011000110101010: color_data = 12'b111011101110;
20'b00100011000110101011: color_data = 12'b111011101110;
20'b00100011000110101100: color_data = 12'b111011101110;
20'b00100011000110101101: color_data = 12'b111011101110;
20'b00100011000110101110: color_data = 12'b111011101110;
20'b00100011000110101111: color_data = 12'b111011101110;
20'b00100011000110110000: color_data = 12'b111011101110;
20'b00100011000110110001: color_data = 12'b111011101110;
20'b00100011000110110010: color_data = 12'b111011101110;
20'b00100011010010010110: color_data = 12'b111011101110;
20'b00100011010010010111: color_data = 12'b111011101110;
20'b00100011010010011000: color_data = 12'b111011101110;
20'b00100011010010011001: color_data = 12'b111011101110;
20'b00100011010010011010: color_data = 12'b111011101110;
20'b00100011010010011011: color_data = 12'b111011101110;
20'b00100011010010011100: color_data = 12'b111011101110;
20'b00100011010010011101: color_data = 12'b111011101110;
20'b00100011010010011110: color_data = 12'b111011101110;
20'b00100011010010011111: color_data = 12'b111011101110;
20'b00100011010010100001: color_data = 12'b111011101110;
20'b00100011010010100010: color_data = 12'b111011101110;
20'b00100011010010100011: color_data = 12'b111011101110;
20'b00100011010010100100: color_data = 12'b111011101110;
20'b00100011010010100101: color_data = 12'b111011101110;
20'b00100011010010100110: color_data = 12'b111011101110;
20'b00100011010010100111: color_data = 12'b111011101110;
20'b00100011010010101000: color_data = 12'b111011101110;
20'b00100011010010101001: color_data = 12'b111011101110;
20'b00100011010010101010: color_data = 12'b111011101110;
20'b00100011010011101110: color_data = 12'b111011101110;
20'b00100011010011101111: color_data = 12'b111011101110;
20'b00100011010011110000: color_data = 12'b111011101110;
20'b00100011010011110001: color_data = 12'b111011101110;
20'b00100011010011110010: color_data = 12'b111011101110;
20'b00100011010011110011: color_data = 12'b111011101110;
20'b00100011010011110100: color_data = 12'b111011101110;
20'b00100011010011110101: color_data = 12'b111011101110;
20'b00100011010011110110: color_data = 12'b111011101110;
20'b00100011010011110111: color_data = 12'b111011101110;
20'b00100011010011111001: color_data = 12'b111011101110;
20'b00100011010011111010: color_data = 12'b111011101110;
20'b00100011010011111011: color_data = 12'b111011101110;
20'b00100011010011111100: color_data = 12'b111011101110;
20'b00100011010011111101: color_data = 12'b111011101110;
20'b00100011010011111110: color_data = 12'b111011101110;
20'b00100011010011111111: color_data = 12'b111011101110;
20'b00100011010100000000: color_data = 12'b111011101110;
20'b00100011010100000001: color_data = 12'b111011101110;
20'b00100011010100000010: color_data = 12'b111011101110;
20'b00100011010100100101: color_data = 12'b111011101110;
20'b00100011010100100110: color_data = 12'b111011101110;
20'b00100011010100100111: color_data = 12'b111011101110;
20'b00100011010100101000: color_data = 12'b111011101110;
20'b00100011010100101001: color_data = 12'b111011101110;
20'b00100011010100101010: color_data = 12'b111011101110;
20'b00100011010100101011: color_data = 12'b111011101110;
20'b00100011010100101100: color_data = 12'b111011101110;
20'b00100011010100101101: color_data = 12'b111011101110;
20'b00100011010100101110: color_data = 12'b111011101110;
20'b00100011010100110000: color_data = 12'b111011101110;
20'b00100011010100110001: color_data = 12'b111011101110;
20'b00100011010100110010: color_data = 12'b111011101110;
20'b00100011010100110011: color_data = 12'b111011101110;
20'b00100011010100110100: color_data = 12'b111011101110;
20'b00100011010100110101: color_data = 12'b111011101110;
20'b00100011010100110110: color_data = 12'b111011101110;
20'b00100011010100110111: color_data = 12'b111011101110;
20'b00100011010100111000: color_data = 12'b111011101110;
20'b00100011010100111001: color_data = 12'b111011101110;
20'b00100011010101000110: color_data = 12'b111011101110;
20'b00100011010101000111: color_data = 12'b111011101110;
20'b00100011010101001000: color_data = 12'b111011101110;
20'b00100011010101001001: color_data = 12'b111011101110;
20'b00100011010101001010: color_data = 12'b111011101110;
20'b00100011010101001011: color_data = 12'b111011101110;
20'b00100011010101001100: color_data = 12'b111011101110;
20'b00100011010101001101: color_data = 12'b111011101110;
20'b00100011010101001110: color_data = 12'b111011101110;
20'b00100011010101001111: color_data = 12'b111011101110;
20'b00100011010101010001: color_data = 12'b111011101110;
20'b00100011010101010010: color_data = 12'b111011101110;
20'b00100011010101010011: color_data = 12'b111011101110;
20'b00100011010101010100: color_data = 12'b111011101110;
20'b00100011010101010101: color_data = 12'b111011101110;
20'b00100011010101010110: color_data = 12'b111011101110;
20'b00100011010101010111: color_data = 12'b111011101110;
20'b00100011010101011000: color_data = 12'b111011101110;
20'b00100011010101011001: color_data = 12'b111011101110;
20'b00100011010101011010: color_data = 12'b111011101110;
20'b00100011010101011100: color_data = 12'b111011101110;
20'b00100011010101011101: color_data = 12'b111011101110;
20'b00100011010101011110: color_data = 12'b111011101110;
20'b00100011010101011111: color_data = 12'b111011101110;
20'b00100011010101100000: color_data = 12'b111011101110;
20'b00100011010101100001: color_data = 12'b111011101110;
20'b00100011010101100010: color_data = 12'b111011101110;
20'b00100011010101100011: color_data = 12'b111011101110;
20'b00100011010101100100: color_data = 12'b111011101110;
20'b00100011010101100101: color_data = 12'b111011101110;
20'b00100011010101100111: color_data = 12'b111011101110;
20'b00100011010101101000: color_data = 12'b111011101110;
20'b00100011010101101001: color_data = 12'b111011101110;
20'b00100011010101101010: color_data = 12'b111011101110;
20'b00100011010101101011: color_data = 12'b111011101110;
20'b00100011010101101100: color_data = 12'b111011101110;
20'b00100011010101101101: color_data = 12'b111011101110;
20'b00100011010101101110: color_data = 12'b111011101110;
20'b00100011010101101111: color_data = 12'b111011101110;
20'b00100011010101110000: color_data = 12'b111011101110;
20'b00100011010101110010: color_data = 12'b111011101110;
20'b00100011010101110011: color_data = 12'b111011101110;
20'b00100011010101110100: color_data = 12'b111011101110;
20'b00100011010101110101: color_data = 12'b111011101110;
20'b00100011010101110110: color_data = 12'b111011101110;
20'b00100011010101110111: color_data = 12'b111011101110;
20'b00100011010101111000: color_data = 12'b111011101110;
20'b00100011010101111001: color_data = 12'b111011101110;
20'b00100011010101111010: color_data = 12'b111011101110;
20'b00100011010101111011: color_data = 12'b111011101110;
20'b00100011010101111101: color_data = 12'b111011101110;
20'b00100011010101111110: color_data = 12'b111011101110;
20'b00100011010101111111: color_data = 12'b111011101110;
20'b00100011010110000000: color_data = 12'b111011101110;
20'b00100011010110000001: color_data = 12'b111011101110;
20'b00100011010110000010: color_data = 12'b111011101110;
20'b00100011010110000011: color_data = 12'b111011101110;
20'b00100011010110000100: color_data = 12'b111011101110;
20'b00100011010110000101: color_data = 12'b111011101110;
20'b00100011010110000110: color_data = 12'b111011101110;
20'b00100011010110001000: color_data = 12'b111011101110;
20'b00100011010110001001: color_data = 12'b111011101110;
20'b00100011010110001010: color_data = 12'b111011101110;
20'b00100011010110001011: color_data = 12'b111011101110;
20'b00100011010110001100: color_data = 12'b111011101110;
20'b00100011010110001101: color_data = 12'b111011101110;
20'b00100011010110001110: color_data = 12'b111011101110;
20'b00100011010110001111: color_data = 12'b111011101110;
20'b00100011010110010000: color_data = 12'b111011101110;
20'b00100011010110010001: color_data = 12'b111011101110;
20'b00100011010110101001: color_data = 12'b111011101110;
20'b00100011010110101010: color_data = 12'b111011101110;
20'b00100011010110101011: color_data = 12'b111011101110;
20'b00100011010110101100: color_data = 12'b111011101110;
20'b00100011010110101101: color_data = 12'b111011101110;
20'b00100011010110101110: color_data = 12'b111011101110;
20'b00100011010110101111: color_data = 12'b111011101110;
20'b00100011010110110000: color_data = 12'b111011101110;
20'b00100011010110110001: color_data = 12'b111011101110;
20'b00100011010110110010: color_data = 12'b111011101110;
20'b00100011100010010110: color_data = 12'b111011101110;
20'b00100011100010010111: color_data = 12'b111011101110;
20'b00100011100010011000: color_data = 12'b111011101110;
20'b00100011100010011001: color_data = 12'b111011101110;
20'b00100011100010011010: color_data = 12'b111011101110;
20'b00100011100010011011: color_data = 12'b111011101110;
20'b00100011100010011100: color_data = 12'b111011101110;
20'b00100011100010011101: color_data = 12'b111011101110;
20'b00100011100010011110: color_data = 12'b111011101110;
20'b00100011100010011111: color_data = 12'b111011101110;
20'b00100011100010100001: color_data = 12'b111011101110;
20'b00100011100010100010: color_data = 12'b111011101110;
20'b00100011100010100011: color_data = 12'b111011101110;
20'b00100011100010100100: color_data = 12'b111011101110;
20'b00100011100010100101: color_data = 12'b111011101110;
20'b00100011100010100110: color_data = 12'b111011101110;
20'b00100011100010100111: color_data = 12'b111011101110;
20'b00100011100010101000: color_data = 12'b111011101110;
20'b00100011100010101001: color_data = 12'b111011101110;
20'b00100011100010101010: color_data = 12'b111011101110;
20'b00100011100011101110: color_data = 12'b111011101110;
20'b00100011100011101111: color_data = 12'b111011101110;
20'b00100011100011110000: color_data = 12'b111011101110;
20'b00100011100011110001: color_data = 12'b111011101110;
20'b00100011100011110010: color_data = 12'b111011101110;
20'b00100011100011110011: color_data = 12'b111011101110;
20'b00100011100011110100: color_data = 12'b111011101110;
20'b00100011100011110101: color_data = 12'b111011101110;
20'b00100011100011110110: color_data = 12'b111011101110;
20'b00100011100011110111: color_data = 12'b111011101110;
20'b00100011100011111001: color_data = 12'b111011101110;
20'b00100011100011111010: color_data = 12'b111011101110;
20'b00100011100011111011: color_data = 12'b111011101110;
20'b00100011100011111100: color_data = 12'b111011101110;
20'b00100011100011111101: color_data = 12'b111011101110;
20'b00100011100011111110: color_data = 12'b111011101110;
20'b00100011100011111111: color_data = 12'b111011101110;
20'b00100011100100000000: color_data = 12'b111011101110;
20'b00100011100100000001: color_data = 12'b111011101110;
20'b00100011100100000010: color_data = 12'b111011101110;
20'b00100011100100100101: color_data = 12'b111011101110;
20'b00100011100100100110: color_data = 12'b111011101110;
20'b00100011100100100111: color_data = 12'b111011101110;
20'b00100011100100101000: color_data = 12'b111011101110;
20'b00100011100100101001: color_data = 12'b111011101110;
20'b00100011100100101010: color_data = 12'b111011101110;
20'b00100011100100101011: color_data = 12'b111011101110;
20'b00100011100100101100: color_data = 12'b111011101110;
20'b00100011100100101101: color_data = 12'b111011101110;
20'b00100011100100101110: color_data = 12'b111011101110;
20'b00100011100100110000: color_data = 12'b111011101110;
20'b00100011100100110001: color_data = 12'b111011101110;
20'b00100011100100110010: color_data = 12'b111011101110;
20'b00100011100100110011: color_data = 12'b111011101110;
20'b00100011100100110100: color_data = 12'b111011101110;
20'b00100011100100110101: color_data = 12'b111011101110;
20'b00100011100100110110: color_data = 12'b111011101110;
20'b00100011100100110111: color_data = 12'b111011101110;
20'b00100011100100111000: color_data = 12'b111011101110;
20'b00100011100100111001: color_data = 12'b111011101110;
20'b00100011100101000110: color_data = 12'b111011101110;
20'b00100011100101000111: color_data = 12'b111011101110;
20'b00100011100101001000: color_data = 12'b111011101110;
20'b00100011100101001001: color_data = 12'b111011101110;
20'b00100011100101001010: color_data = 12'b111011101110;
20'b00100011100101001011: color_data = 12'b111011101110;
20'b00100011100101001100: color_data = 12'b111011101110;
20'b00100011100101001101: color_data = 12'b111011101110;
20'b00100011100101001110: color_data = 12'b111011101110;
20'b00100011100101001111: color_data = 12'b111011101110;
20'b00100011100101010001: color_data = 12'b111011101110;
20'b00100011100101010010: color_data = 12'b111011101110;
20'b00100011100101010011: color_data = 12'b111011101110;
20'b00100011100101010100: color_data = 12'b111011101110;
20'b00100011100101010101: color_data = 12'b111011101110;
20'b00100011100101010110: color_data = 12'b111011101110;
20'b00100011100101010111: color_data = 12'b111011101110;
20'b00100011100101011000: color_data = 12'b111011101110;
20'b00100011100101011001: color_data = 12'b111011101110;
20'b00100011100101011010: color_data = 12'b111011101110;
20'b00100011100101011100: color_data = 12'b111011101110;
20'b00100011100101011101: color_data = 12'b111011101110;
20'b00100011100101011110: color_data = 12'b111011101110;
20'b00100011100101011111: color_data = 12'b111011101110;
20'b00100011100101100000: color_data = 12'b111011101110;
20'b00100011100101100001: color_data = 12'b111011101110;
20'b00100011100101100010: color_data = 12'b111011101110;
20'b00100011100101100011: color_data = 12'b111011101110;
20'b00100011100101100100: color_data = 12'b111011101110;
20'b00100011100101100101: color_data = 12'b111011101110;
20'b00100011100101100111: color_data = 12'b111011101110;
20'b00100011100101101000: color_data = 12'b111011101110;
20'b00100011100101101001: color_data = 12'b111011101110;
20'b00100011100101101010: color_data = 12'b111011101110;
20'b00100011100101101011: color_data = 12'b111011101110;
20'b00100011100101101100: color_data = 12'b111011101110;
20'b00100011100101101101: color_data = 12'b111011101110;
20'b00100011100101101110: color_data = 12'b111011101110;
20'b00100011100101101111: color_data = 12'b111011101110;
20'b00100011100101110000: color_data = 12'b111011101110;
20'b00100011100101110010: color_data = 12'b111011101110;
20'b00100011100101110011: color_data = 12'b111011101110;
20'b00100011100101110100: color_data = 12'b111011101110;
20'b00100011100101110101: color_data = 12'b111011101110;
20'b00100011100101110110: color_data = 12'b111011101110;
20'b00100011100101110111: color_data = 12'b111011101110;
20'b00100011100101111000: color_data = 12'b111011101110;
20'b00100011100101111001: color_data = 12'b111011101110;
20'b00100011100101111010: color_data = 12'b111011101110;
20'b00100011100101111011: color_data = 12'b111011101110;
20'b00100011100101111101: color_data = 12'b111011101110;
20'b00100011100101111110: color_data = 12'b111011101110;
20'b00100011100101111111: color_data = 12'b111011101110;
20'b00100011100110000000: color_data = 12'b111011101110;
20'b00100011100110000001: color_data = 12'b111011101110;
20'b00100011100110000010: color_data = 12'b111011101110;
20'b00100011100110000011: color_data = 12'b111011101110;
20'b00100011100110000100: color_data = 12'b111011101110;
20'b00100011100110000101: color_data = 12'b111011101110;
20'b00100011100110000110: color_data = 12'b111011101110;
20'b00100011100110001000: color_data = 12'b111011101110;
20'b00100011100110001001: color_data = 12'b111011101110;
20'b00100011100110001010: color_data = 12'b111011101110;
20'b00100011100110001011: color_data = 12'b111011101110;
20'b00100011100110001100: color_data = 12'b111011101110;
20'b00100011100110001101: color_data = 12'b111011101110;
20'b00100011100110001110: color_data = 12'b111011101110;
20'b00100011100110001111: color_data = 12'b111011101110;
20'b00100011100110010000: color_data = 12'b111011101110;
20'b00100011100110010001: color_data = 12'b111011101110;
20'b00100011100110101001: color_data = 12'b111011101110;
20'b00100011100110101010: color_data = 12'b111011101110;
20'b00100011100110101011: color_data = 12'b111011101110;
20'b00100011100110101100: color_data = 12'b111011101110;
20'b00100011100110101101: color_data = 12'b111011101110;
20'b00100011100110101110: color_data = 12'b111011101110;
20'b00100011100110101111: color_data = 12'b111011101110;
20'b00100011100110110000: color_data = 12'b111011101110;
20'b00100011100110110001: color_data = 12'b111011101110;
20'b00100011100110110010: color_data = 12'b111011101110;
20'b00100011110010010110: color_data = 12'b111011101110;
20'b00100011110010010111: color_data = 12'b111011101110;
20'b00100011110010011000: color_data = 12'b111011101110;
20'b00100011110010011001: color_data = 12'b111011101110;
20'b00100011110010011010: color_data = 12'b111011101110;
20'b00100011110010011011: color_data = 12'b111011101110;
20'b00100011110010011100: color_data = 12'b111011101110;
20'b00100011110010011101: color_data = 12'b111011101110;
20'b00100011110010011110: color_data = 12'b111011101110;
20'b00100011110010011111: color_data = 12'b111011101110;
20'b00100011110010100001: color_data = 12'b111011101110;
20'b00100011110010100010: color_data = 12'b111011101110;
20'b00100011110010100011: color_data = 12'b111011101110;
20'b00100011110010100100: color_data = 12'b111011101110;
20'b00100011110010100101: color_data = 12'b111011101110;
20'b00100011110010100110: color_data = 12'b111011101110;
20'b00100011110010100111: color_data = 12'b111011101110;
20'b00100011110010101000: color_data = 12'b111011101110;
20'b00100011110010101001: color_data = 12'b111011101110;
20'b00100011110010101010: color_data = 12'b111011101110;
20'b00100011110011101110: color_data = 12'b111011101110;
20'b00100011110011101111: color_data = 12'b111011101110;
20'b00100011110011110000: color_data = 12'b111011101110;
20'b00100011110011110001: color_data = 12'b111011101110;
20'b00100011110011110010: color_data = 12'b111011101110;
20'b00100011110011110011: color_data = 12'b111011101110;
20'b00100011110011110100: color_data = 12'b111011101110;
20'b00100011110011110101: color_data = 12'b111011101110;
20'b00100011110011110110: color_data = 12'b111011101110;
20'b00100011110011110111: color_data = 12'b111011101110;
20'b00100011110011111001: color_data = 12'b111011101110;
20'b00100011110011111010: color_data = 12'b111011101110;
20'b00100011110011111011: color_data = 12'b111011101110;
20'b00100011110011111100: color_data = 12'b111011101110;
20'b00100011110011111101: color_data = 12'b111011101110;
20'b00100011110011111110: color_data = 12'b111011101110;
20'b00100011110011111111: color_data = 12'b111011101110;
20'b00100011110100000000: color_data = 12'b111011101110;
20'b00100011110100000001: color_data = 12'b111011101110;
20'b00100011110100000010: color_data = 12'b111011101110;
20'b00100011110100100101: color_data = 12'b111011101110;
20'b00100011110100100110: color_data = 12'b111011101110;
20'b00100011110100100111: color_data = 12'b111011101110;
20'b00100011110100101000: color_data = 12'b111011101110;
20'b00100011110100101001: color_data = 12'b111011101110;
20'b00100011110100101010: color_data = 12'b111011101110;
20'b00100011110100101011: color_data = 12'b111011101110;
20'b00100011110100101100: color_data = 12'b111011101110;
20'b00100011110100101101: color_data = 12'b111011101110;
20'b00100011110100101110: color_data = 12'b111011101110;
20'b00100011110100110000: color_data = 12'b111011101110;
20'b00100011110100110001: color_data = 12'b111011101110;
20'b00100011110100110010: color_data = 12'b111011101110;
20'b00100011110100110011: color_data = 12'b111011101110;
20'b00100011110100110100: color_data = 12'b111011101110;
20'b00100011110100110101: color_data = 12'b111011101110;
20'b00100011110100110110: color_data = 12'b111011101110;
20'b00100011110100110111: color_data = 12'b111011101110;
20'b00100011110100111000: color_data = 12'b111011101110;
20'b00100011110100111001: color_data = 12'b111011101110;
20'b00100011110101000110: color_data = 12'b111011101110;
20'b00100011110101000111: color_data = 12'b111011101110;
20'b00100011110101001000: color_data = 12'b111011101110;
20'b00100011110101001001: color_data = 12'b111011101110;
20'b00100011110101001010: color_data = 12'b111011101110;
20'b00100011110101001011: color_data = 12'b111011101110;
20'b00100011110101001100: color_data = 12'b111011101110;
20'b00100011110101001101: color_data = 12'b111011101110;
20'b00100011110101001110: color_data = 12'b111011101110;
20'b00100011110101001111: color_data = 12'b111011101110;
20'b00100011110101010001: color_data = 12'b111011101110;
20'b00100011110101010010: color_data = 12'b111011101110;
20'b00100011110101010011: color_data = 12'b111011101110;
20'b00100011110101010100: color_data = 12'b111011101110;
20'b00100011110101010101: color_data = 12'b111011101110;
20'b00100011110101010110: color_data = 12'b111011101110;
20'b00100011110101010111: color_data = 12'b111011101110;
20'b00100011110101011000: color_data = 12'b111011101110;
20'b00100011110101011001: color_data = 12'b111011101110;
20'b00100011110101011010: color_data = 12'b111011101110;
20'b00100011110101011100: color_data = 12'b111011101110;
20'b00100011110101011101: color_data = 12'b111011101110;
20'b00100011110101011110: color_data = 12'b111011101110;
20'b00100011110101011111: color_data = 12'b111011101110;
20'b00100011110101100000: color_data = 12'b111011101110;
20'b00100011110101100001: color_data = 12'b111011101110;
20'b00100011110101100010: color_data = 12'b111011101110;
20'b00100011110101100011: color_data = 12'b111011101110;
20'b00100011110101100100: color_data = 12'b111011101110;
20'b00100011110101100101: color_data = 12'b111011101110;
20'b00100011110101100111: color_data = 12'b111011101110;
20'b00100011110101101000: color_data = 12'b111011101110;
20'b00100011110101101001: color_data = 12'b111011101110;
20'b00100011110101101010: color_data = 12'b111011101110;
20'b00100011110101101011: color_data = 12'b111011101110;
20'b00100011110101101100: color_data = 12'b111011101110;
20'b00100011110101101101: color_data = 12'b111011101110;
20'b00100011110101101110: color_data = 12'b111011101110;
20'b00100011110101101111: color_data = 12'b111011101110;
20'b00100011110101110000: color_data = 12'b111011101110;
20'b00100011110101110010: color_data = 12'b111011101110;
20'b00100011110101110011: color_data = 12'b111011101110;
20'b00100011110101110100: color_data = 12'b111011101110;
20'b00100011110101110101: color_data = 12'b111011101110;
20'b00100011110101110110: color_data = 12'b111011101110;
20'b00100011110101110111: color_data = 12'b111011101110;
20'b00100011110101111000: color_data = 12'b111011101110;
20'b00100011110101111001: color_data = 12'b111011101110;
20'b00100011110101111010: color_data = 12'b111011101110;
20'b00100011110101111011: color_data = 12'b111011101110;
20'b00100011110101111101: color_data = 12'b111011101110;
20'b00100011110101111110: color_data = 12'b111011101110;
20'b00100011110101111111: color_data = 12'b111011101110;
20'b00100011110110000000: color_data = 12'b111011101110;
20'b00100011110110000001: color_data = 12'b111011101110;
20'b00100011110110000010: color_data = 12'b111011101110;
20'b00100011110110000011: color_data = 12'b111011101110;
20'b00100011110110000100: color_data = 12'b111011101110;
20'b00100011110110000101: color_data = 12'b111011101110;
20'b00100011110110000110: color_data = 12'b111011101110;
20'b00100011110110001000: color_data = 12'b111011101110;
20'b00100011110110001001: color_data = 12'b111011101110;
20'b00100011110110001010: color_data = 12'b111011101110;
20'b00100011110110001011: color_data = 12'b111011101110;
20'b00100011110110001100: color_data = 12'b111011101110;
20'b00100011110110001101: color_data = 12'b111011101110;
20'b00100011110110001110: color_data = 12'b111011101110;
20'b00100011110110001111: color_data = 12'b111011101110;
20'b00100011110110010000: color_data = 12'b111011101110;
20'b00100011110110010001: color_data = 12'b111011101110;
20'b00100011110110101001: color_data = 12'b111011101110;
20'b00100011110110101010: color_data = 12'b111011101110;
20'b00100011110110101011: color_data = 12'b111011101110;
20'b00100011110110101100: color_data = 12'b111011101110;
20'b00100011110110101101: color_data = 12'b111011101110;
20'b00100011110110101110: color_data = 12'b111011101110;
20'b00100011110110101111: color_data = 12'b111011101110;
20'b00100011110110110000: color_data = 12'b111011101110;
20'b00100011110110110001: color_data = 12'b111011101110;
20'b00100011110110110010: color_data = 12'b111011101110;
20'b00100100000010010110: color_data = 12'b111011101110;
20'b00100100000010010111: color_data = 12'b111011101110;
20'b00100100000010011000: color_data = 12'b111011101110;
20'b00100100000010011001: color_data = 12'b111011101110;
20'b00100100000010011010: color_data = 12'b111011101110;
20'b00100100000010011011: color_data = 12'b111011101110;
20'b00100100000010011100: color_data = 12'b111011101110;
20'b00100100000010011101: color_data = 12'b111011101110;
20'b00100100000010011110: color_data = 12'b111011101110;
20'b00100100000010011111: color_data = 12'b111011101110;
20'b00100100000010100001: color_data = 12'b111011101110;
20'b00100100000010100010: color_data = 12'b111011101110;
20'b00100100000010100011: color_data = 12'b111011101110;
20'b00100100000010100100: color_data = 12'b111011101110;
20'b00100100000010100101: color_data = 12'b111011101110;
20'b00100100000010100110: color_data = 12'b111011101110;
20'b00100100000010100111: color_data = 12'b111011101110;
20'b00100100000010101000: color_data = 12'b111011101110;
20'b00100100000010101001: color_data = 12'b111011101110;
20'b00100100000010101010: color_data = 12'b111011101110;
20'b00100100000011101110: color_data = 12'b111011101110;
20'b00100100000011101111: color_data = 12'b111011101110;
20'b00100100000011110000: color_data = 12'b111011101110;
20'b00100100000011110001: color_data = 12'b111011101110;
20'b00100100000011110010: color_data = 12'b111011101110;
20'b00100100000011110011: color_data = 12'b111011101110;
20'b00100100000011110100: color_data = 12'b111011101110;
20'b00100100000011110101: color_data = 12'b111011101110;
20'b00100100000011110110: color_data = 12'b111011101110;
20'b00100100000011110111: color_data = 12'b111011101110;
20'b00100100000011111001: color_data = 12'b111011101110;
20'b00100100000011111010: color_data = 12'b111011101110;
20'b00100100000011111011: color_data = 12'b111011101110;
20'b00100100000011111100: color_data = 12'b111011101110;
20'b00100100000011111101: color_data = 12'b111011101110;
20'b00100100000011111110: color_data = 12'b111011101110;
20'b00100100000011111111: color_data = 12'b111011101110;
20'b00100100000100000000: color_data = 12'b111011101110;
20'b00100100000100000001: color_data = 12'b111011101110;
20'b00100100000100000010: color_data = 12'b111011101110;
20'b00100100000100100101: color_data = 12'b111011101110;
20'b00100100000100100110: color_data = 12'b111011101110;
20'b00100100000100100111: color_data = 12'b111011101110;
20'b00100100000100101000: color_data = 12'b111011101110;
20'b00100100000100101001: color_data = 12'b111011101110;
20'b00100100000100101010: color_data = 12'b111011101110;
20'b00100100000100101011: color_data = 12'b111011101110;
20'b00100100000100101100: color_data = 12'b111011101110;
20'b00100100000100101101: color_data = 12'b111011101110;
20'b00100100000100101110: color_data = 12'b111011101110;
20'b00100100000100110000: color_data = 12'b111011101110;
20'b00100100000100110001: color_data = 12'b111011101110;
20'b00100100000100110010: color_data = 12'b111011101110;
20'b00100100000100110011: color_data = 12'b111011101110;
20'b00100100000100110100: color_data = 12'b111011101110;
20'b00100100000100110101: color_data = 12'b111011101110;
20'b00100100000100110110: color_data = 12'b111011101110;
20'b00100100000100110111: color_data = 12'b111011101110;
20'b00100100000100111000: color_data = 12'b111011101110;
20'b00100100000100111001: color_data = 12'b111011101110;
20'b00100100000101000110: color_data = 12'b111011101110;
20'b00100100000101000111: color_data = 12'b111011101110;
20'b00100100000101001000: color_data = 12'b111011101110;
20'b00100100000101001001: color_data = 12'b111011101110;
20'b00100100000101001010: color_data = 12'b111011101110;
20'b00100100000101001011: color_data = 12'b111011101110;
20'b00100100000101001100: color_data = 12'b111011101110;
20'b00100100000101001101: color_data = 12'b111011101110;
20'b00100100000101001110: color_data = 12'b111011101110;
20'b00100100000101001111: color_data = 12'b111011101110;
20'b00100100000101010001: color_data = 12'b111011101110;
20'b00100100000101010010: color_data = 12'b111011101110;
20'b00100100000101010011: color_data = 12'b111011101110;
20'b00100100000101010100: color_data = 12'b111011101110;
20'b00100100000101010101: color_data = 12'b111011101110;
20'b00100100000101010110: color_data = 12'b111011101110;
20'b00100100000101010111: color_data = 12'b111011101110;
20'b00100100000101011000: color_data = 12'b111011101110;
20'b00100100000101011001: color_data = 12'b111011101110;
20'b00100100000101011010: color_data = 12'b111011101110;
20'b00100100000101011100: color_data = 12'b111011101110;
20'b00100100000101011101: color_data = 12'b111011101110;
20'b00100100000101011110: color_data = 12'b111011101110;
20'b00100100000101011111: color_data = 12'b111011101110;
20'b00100100000101100000: color_data = 12'b111011101110;
20'b00100100000101100001: color_data = 12'b111011101110;
20'b00100100000101100010: color_data = 12'b111011101110;
20'b00100100000101100011: color_data = 12'b111011101110;
20'b00100100000101100100: color_data = 12'b111011101110;
20'b00100100000101100101: color_data = 12'b111011101110;
20'b00100100000101100111: color_data = 12'b111011101110;
20'b00100100000101101000: color_data = 12'b111011101110;
20'b00100100000101101001: color_data = 12'b111011101110;
20'b00100100000101101010: color_data = 12'b111011101110;
20'b00100100000101101011: color_data = 12'b111011101110;
20'b00100100000101101100: color_data = 12'b111011101110;
20'b00100100000101101101: color_data = 12'b111011101110;
20'b00100100000101101110: color_data = 12'b111011101110;
20'b00100100000101101111: color_data = 12'b111011101110;
20'b00100100000101110000: color_data = 12'b111011101110;
20'b00100100000101110010: color_data = 12'b111011101110;
20'b00100100000101110011: color_data = 12'b111011101110;
20'b00100100000101110100: color_data = 12'b111011101110;
20'b00100100000101110101: color_data = 12'b111011101110;
20'b00100100000101110110: color_data = 12'b111011101110;
20'b00100100000101110111: color_data = 12'b111011101110;
20'b00100100000101111000: color_data = 12'b111011101110;
20'b00100100000101111001: color_data = 12'b111011101110;
20'b00100100000101111010: color_data = 12'b111011101110;
20'b00100100000101111011: color_data = 12'b111011101110;
20'b00100100000101111101: color_data = 12'b111011101110;
20'b00100100000101111110: color_data = 12'b111011101110;
20'b00100100000101111111: color_data = 12'b111011101110;
20'b00100100000110000000: color_data = 12'b111011101110;
20'b00100100000110000001: color_data = 12'b111011101110;
20'b00100100000110000010: color_data = 12'b111011101110;
20'b00100100000110000011: color_data = 12'b111011101110;
20'b00100100000110000100: color_data = 12'b111011101110;
20'b00100100000110000101: color_data = 12'b111011101110;
20'b00100100000110000110: color_data = 12'b111011101110;
20'b00100100000110001000: color_data = 12'b111011101110;
20'b00100100000110001001: color_data = 12'b111011101110;
20'b00100100000110001010: color_data = 12'b111011101110;
20'b00100100000110001011: color_data = 12'b111011101110;
20'b00100100000110001100: color_data = 12'b111011101110;
20'b00100100000110001101: color_data = 12'b111011101110;
20'b00100100000110001110: color_data = 12'b111011101110;
20'b00100100000110001111: color_data = 12'b111011101110;
20'b00100100000110010000: color_data = 12'b111011101110;
20'b00100100000110010001: color_data = 12'b111011101110;
20'b00100100000110101001: color_data = 12'b111011101110;
20'b00100100000110101010: color_data = 12'b111011101110;
20'b00100100000110101011: color_data = 12'b111011101110;
20'b00100100000110101100: color_data = 12'b111011101110;
20'b00100100000110101101: color_data = 12'b111011101110;
20'b00100100000110101110: color_data = 12'b111011101110;
20'b00100100000110101111: color_data = 12'b111011101110;
20'b00100100000110110000: color_data = 12'b111011101110;
20'b00100100000110110001: color_data = 12'b111011101110;
20'b00100100000110110010: color_data = 12'b111011101110;
20'b00100100010010010110: color_data = 12'b111011101110;
20'b00100100010010010111: color_data = 12'b111011101110;
20'b00100100010010011000: color_data = 12'b111011101110;
20'b00100100010010011001: color_data = 12'b111011101110;
20'b00100100010010011010: color_data = 12'b111011101110;
20'b00100100010010011011: color_data = 12'b111011101110;
20'b00100100010010011100: color_data = 12'b111011101110;
20'b00100100010010011101: color_data = 12'b111011101110;
20'b00100100010010011110: color_data = 12'b111011101110;
20'b00100100010010011111: color_data = 12'b111011101110;
20'b00100100010010100001: color_data = 12'b111011101110;
20'b00100100010010100010: color_data = 12'b111011101110;
20'b00100100010010100011: color_data = 12'b111011101110;
20'b00100100010010100100: color_data = 12'b111011101110;
20'b00100100010010100101: color_data = 12'b111011101110;
20'b00100100010010100110: color_data = 12'b111011101110;
20'b00100100010010100111: color_data = 12'b111011101110;
20'b00100100010010101000: color_data = 12'b111011101110;
20'b00100100010010101001: color_data = 12'b111011101110;
20'b00100100010010101010: color_data = 12'b111011101110;
20'b00100100010011101110: color_data = 12'b111011101110;
20'b00100100010011101111: color_data = 12'b111011101110;
20'b00100100010011110000: color_data = 12'b111011101110;
20'b00100100010011110001: color_data = 12'b111011101110;
20'b00100100010011110010: color_data = 12'b111011101110;
20'b00100100010011110011: color_data = 12'b111011101110;
20'b00100100010011110100: color_data = 12'b111011101110;
20'b00100100010011110101: color_data = 12'b111011101110;
20'b00100100010011110110: color_data = 12'b111011101110;
20'b00100100010011110111: color_data = 12'b111011101110;
20'b00100100010011111001: color_data = 12'b111011101110;
20'b00100100010011111010: color_data = 12'b111011101110;
20'b00100100010011111011: color_data = 12'b111011101110;
20'b00100100010011111100: color_data = 12'b111011101110;
20'b00100100010011111101: color_data = 12'b111011101110;
20'b00100100010011111110: color_data = 12'b111011101110;
20'b00100100010011111111: color_data = 12'b111011101110;
20'b00100100010100000000: color_data = 12'b111011101110;
20'b00100100010100000001: color_data = 12'b111011101110;
20'b00100100010100000010: color_data = 12'b111011101110;
20'b00100100010100100101: color_data = 12'b111011101110;
20'b00100100010100100110: color_data = 12'b111011101110;
20'b00100100010100100111: color_data = 12'b111011101110;
20'b00100100010100101000: color_data = 12'b111011101110;
20'b00100100010100101001: color_data = 12'b111011101110;
20'b00100100010100101010: color_data = 12'b111011101110;
20'b00100100010100101011: color_data = 12'b111011101110;
20'b00100100010100101100: color_data = 12'b111011101110;
20'b00100100010100101101: color_data = 12'b111011101110;
20'b00100100010100101110: color_data = 12'b111011101110;
20'b00100100010100110000: color_data = 12'b111011101110;
20'b00100100010100110001: color_data = 12'b111011101110;
20'b00100100010100110010: color_data = 12'b111011101110;
20'b00100100010100110011: color_data = 12'b111011101110;
20'b00100100010100110100: color_data = 12'b111011101110;
20'b00100100010100110101: color_data = 12'b111011101110;
20'b00100100010100110110: color_data = 12'b111011101110;
20'b00100100010100110111: color_data = 12'b111011101110;
20'b00100100010100111000: color_data = 12'b111011101110;
20'b00100100010100111001: color_data = 12'b111011101110;
20'b00100100010101000110: color_data = 12'b111011101110;
20'b00100100010101000111: color_data = 12'b111011101110;
20'b00100100010101001000: color_data = 12'b111011101110;
20'b00100100010101001001: color_data = 12'b111011101110;
20'b00100100010101001010: color_data = 12'b111011101110;
20'b00100100010101001011: color_data = 12'b111011101110;
20'b00100100010101001100: color_data = 12'b111011101110;
20'b00100100010101001101: color_data = 12'b111011101110;
20'b00100100010101001110: color_data = 12'b111011101110;
20'b00100100010101001111: color_data = 12'b111011101110;
20'b00100100010101010001: color_data = 12'b111011101110;
20'b00100100010101010010: color_data = 12'b111011101110;
20'b00100100010101010011: color_data = 12'b111011101110;
20'b00100100010101010100: color_data = 12'b111011101110;
20'b00100100010101010101: color_data = 12'b111011101110;
20'b00100100010101010110: color_data = 12'b111011101110;
20'b00100100010101010111: color_data = 12'b111011101110;
20'b00100100010101011000: color_data = 12'b111011101110;
20'b00100100010101011001: color_data = 12'b111011101110;
20'b00100100010101011010: color_data = 12'b111011101110;
20'b00100100010101011100: color_data = 12'b111011101110;
20'b00100100010101011101: color_data = 12'b111011101110;
20'b00100100010101011110: color_data = 12'b111011101110;
20'b00100100010101011111: color_data = 12'b111011101110;
20'b00100100010101100000: color_data = 12'b111011101110;
20'b00100100010101100001: color_data = 12'b111011101110;
20'b00100100010101100010: color_data = 12'b111011101110;
20'b00100100010101100011: color_data = 12'b111011101110;
20'b00100100010101100100: color_data = 12'b111011101110;
20'b00100100010101100101: color_data = 12'b111011101110;
20'b00100100010101100111: color_data = 12'b111011101110;
20'b00100100010101101000: color_data = 12'b111011101110;
20'b00100100010101101001: color_data = 12'b111011101110;
20'b00100100010101101010: color_data = 12'b111011101110;
20'b00100100010101101011: color_data = 12'b111011101110;
20'b00100100010101101100: color_data = 12'b111011101110;
20'b00100100010101101101: color_data = 12'b111011101110;
20'b00100100010101101110: color_data = 12'b111011101110;
20'b00100100010101101111: color_data = 12'b111011101110;
20'b00100100010101110000: color_data = 12'b111011101110;
20'b00100100010101110010: color_data = 12'b111011101110;
20'b00100100010101110011: color_data = 12'b111011101110;
20'b00100100010101110100: color_data = 12'b111011101110;
20'b00100100010101110101: color_data = 12'b111011101110;
20'b00100100010101110110: color_data = 12'b111011101110;
20'b00100100010101110111: color_data = 12'b111011101110;
20'b00100100010101111000: color_data = 12'b111011101110;
20'b00100100010101111001: color_data = 12'b111011101110;
20'b00100100010101111010: color_data = 12'b111011101110;
20'b00100100010101111011: color_data = 12'b111011101110;
20'b00100100010101111101: color_data = 12'b111011101110;
20'b00100100010101111110: color_data = 12'b111011101110;
20'b00100100010101111111: color_data = 12'b111011101110;
20'b00100100010110000000: color_data = 12'b111011101110;
20'b00100100010110000001: color_data = 12'b111011101110;
20'b00100100010110000010: color_data = 12'b111011101110;
20'b00100100010110000011: color_data = 12'b111011101110;
20'b00100100010110000100: color_data = 12'b111011101110;
20'b00100100010110000101: color_data = 12'b111011101110;
20'b00100100010110000110: color_data = 12'b111011101110;
20'b00100100010110001000: color_data = 12'b111011101110;
20'b00100100010110001001: color_data = 12'b111011101110;
20'b00100100010110001010: color_data = 12'b111011101110;
20'b00100100010110001011: color_data = 12'b111011101110;
20'b00100100010110001100: color_data = 12'b111011101110;
20'b00100100010110001101: color_data = 12'b111011101110;
20'b00100100010110001110: color_data = 12'b111011101110;
20'b00100100010110001111: color_data = 12'b111011101110;
20'b00100100010110010000: color_data = 12'b111011101110;
20'b00100100010110010001: color_data = 12'b111011101110;
20'b00100100010110101001: color_data = 12'b111011101110;
20'b00100100010110101010: color_data = 12'b111011101110;
20'b00100100010110101011: color_data = 12'b111011101110;
20'b00100100010110101100: color_data = 12'b111011101110;
20'b00100100010110101101: color_data = 12'b111011101110;
20'b00100100010110101110: color_data = 12'b111011101110;
20'b00100100010110101111: color_data = 12'b111011101110;
20'b00100100010110110000: color_data = 12'b111011101110;
20'b00100100010110110001: color_data = 12'b111011101110;
20'b00100100010110110010: color_data = 12'b111011101110;
20'b00100100110010010110: color_data = 12'b111011101110;
20'b00100100110010010111: color_data = 12'b111011101110;
20'b00100100110010011000: color_data = 12'b111011101110;
20'b00100100110010011001: color_data = 12'b111011101110;
20'b00100100110010011010: color_data = 12'b111011101110;
20'b00100100110010011011: color_data = 12'b111011101110;
20'b00100100110010011100: color_data = 12'b111011101110;
20'b00100100110010011101: color_data = 12'b111011101110;
20'b00100100110010011110: color_data = 12'b111011101110;
20'b00100100110010011111: color_data = 12'b111011101110;
20'b00100100110010100001: color_data = 12'b111011101110;
20'b00100100110010100010: color_data = 12'b111011101110;
20'b00100100110010100011: color_data = 12'b111011101110;
20'b00100100110010100100: color_data = 12'b111011101110;
20'b00100100110010100101: color_data = 12'b111011101110;
20'b00100100110010100110: color_data = 12'b111011101110;
20'b00100100110010100111: color_data = 12'b111011101110;
20'b00100100110010101000: color_data = 12'b111011101110;
20'b00100100110010101001: color_data = 12'b111011101110;
20'b00100100110010101010: color_data = 12'b111011101110;
20'b00100100110011101110: color_data = 12'b111011101110;
20'b00100100110011101111: color_data = 12'b111011101110;
20'b00100100110011110000: color_data = 12'b111011101110;
20'b00100100110011110001: color_data = 12'b111011101110;
20'b00100100110011110010: color_data = 12'b111011101110;
20'b00100100110011110011: color_data = 12'b111011101110;
20'b00100100110011110100: color_data = 12'b111011101110;
20'b00100100110011110101: color_data = 12'b111011101110;
20'b00100100110011110110: color_data = 12'b111011101110;
20'b00100100110011110111: color_data = 12'b111011101110;
20'b00100100110011111001: color_data = 12'b111011101110;
20'b00100100110011111010: color_data = 12'b111011101110;
20'b00100100110011111011: color_data = 12'b111011101110;
20'b00100100110011111100: color_data = 12'b111011101110;
20'b00100100110011111101: color_data = 12'b111011101110;
20'b00100100110011111110: color_data = 12'b111011101110;
20'b00100100110011111111: color_data = 12'b111011101110;
20'b00100100110100000000: color_data = 12'b111011101110;
20'b00100100110100000001: color_data = 12'b111011101110;
20'b00100100110100000010: color_data = 12'b111011101110;
20'b00100100110100100101: color_data = 12'b111011101110;
20'b00100100110100100110: color_data = 12'b111011101110;
20'b00100100110100100111: color_data = 12'b111011101110;
20'b00100100110100101000: color_data = 12'b111011101110;
20'b00100100110100101001: color_data = 12'b111011101110;
20'b00100100110100101010: color_data = 12'b111011101110;
20'b00100100110100101011: color_data = 12'b111011101110;
20'b00100100110100101100: color_data = 12'b111011101110;
20'b00100100110100101101: color_data = 12'b111011101110;
20'b00100100110100101110: color_data = 12'b111011101110;
20'b00100100110100110000: color_data = 12'b111011101110;
20'b00100100110100110001: color_data = 12'b111011101110;
20'b00100100110100110010: color_data = 12'b111011101110;
20'b00100100110100110011: color_data = 12'b111011101110;
20'b00100100110100110100: color_data = 12'b111011101110;
20'b00100100110100110101: color_data = 12'b111011101110;
20'b00100100110100110110: color_data = 12'b111011101110;
20'b00100100110100110111: color_data = 12'b111011101110;
20'b00100100110100111000: color_data = 12'b111011101110;
20'b00100100110100111001: color_data = 12'b111011101110;
20'b00100100110101000110: color_data = 12'b111011101110;
20'b00100100110101000111: color_data = 12'b111011101110;
20'b00100100110101001000: color_data = 12'b111011101110;
20'b00100100110101001001: color_data = 12'b111011101110;
20'b00100100110101001010: color_data = 12'b111011101110;
20'b00100100110101001011: color_data = 12'b111011101110;
20'b00100100110101001100: color_data = 12'b111011101110;
20'b00100100110101001101: color_data = 12'b111011101110;
20'b00100100110101001110: color_data = 12'b111011101110;
20'b00100100110101001111: color_data = 12'b111011101110;
20'b00100100110101010001: color_data = 12'b111011101110;
20'b00100100110101010010: color_data = 12'b111011101110;
20'b00100100110101010011: color_data = 12'b111011101110;
20'b00100100110101010100: color_data = 12'b111011101110;
20'b00100100110101010101: color_data = 12'b111011101110;
20'b00100100110101010110: color_data = 12'b111011101110;
20'b00100100110101010111: color_data = 12'b111011101110;
20'b00100100110101011000: color_data = 12'b111011101110;
20'b00100100110101011001: color_data = 12'b111011101110;
20'b00100100110101011010: color_data = 12'b111011101110;
20'b00100100110101100111: color_data = 12'b111011101110;
20'b00100100110101101000: color_data = 12'b111011101110;
20'b00100100110101101001: color_data = 12'b111011101110;
20'b00100100110101101010: color_data = 12'b111011101110;
20'b00100100110101101011: color_data = 12'b111011101110;
20'b00100100110101101100: color_data = 12'b111011101110;
20'b00100100110101101101: color_data = 12'b111011101110;
20'b00100100110101101110: color_data = 12'b111011101110;
20'b00100100110101101111: color_data = 12'b111011101110;
20'b00100100110101110000: color_data = 12'b111011101110;
20'b00100100110101111101: color_data = 12'b111011101110;
20'b00100100110101111110: color_data = 12'b111011101110;
20'b00100100110101111111: color_data = 12'b111011101110;
20'b00100100110110000000: color_data = 12'b111011101110;
20'b00100100110110000001: color_data = 12'b111011101110;
20'b00100100110110000010: color_data = 12'b111011101110;
20'b00100100110110000011: color_data = 12'b111011101110;
20'b00100100110110000100: color_data = 12'b111011101110;
20'b00100100110110000101: color_data = 12'b111011101110;
20'b00100100110110000110: color_data = 12'b111011101110;
20'b00100100110110001000: color_data = 12'b111011101110;
20'b00100100110110001001: color_data = 12'b111011101110;
20'b00100100110110001010: color_data = 12'b111011101110;
20'b00100100110110001011: color_data = 12'b111011101110;
20'b00100100110110001100: color_data = 12'b111011101110;
20'b00100100110110001101: color_data = 12'b111011101110;
20'b00100100110110001110: color_data = 12'b111011101110;
20'b00100100110110001111: color_data = 12'b111011101110;
20'b00100100110110010000: color_data = 12'b111011101110;
20'b00100100110110010001: color_data = 12'b111011101110;
20'b00100100110110011110: color_data = 12'b111011101110;
20'b00100100110110011111: color_data = 12'b111011101110;
20'b00100100110110100000: color_data = 12'b111011101110;
20'b00100100110110100001: color_data = 12'b111011101110;
20'b00100100110110100010: color_data = 12'b111011101110;
20'b00100100110110100011: color_data = 12'b111011101110;
20'b00100100110110100100: color_data = 12'b111011101110;
20'b00100100110110100101: color_data = 12'b111011101110;
20'b00100100110110100110: color_data = 12'b111011101110;
20'b00100100110110100111: color_data = 12'b111011101110;
20'b00100100110110101001: color_data = 12'b111011101110;
20'b00100100110110101010: color_data = 12'b111011101110;
20'b00100100110110101011: color_data = 12'b111011101110;
20'b00100100110110101100: color_data = 12'b111011101110;
20'b00100100110110101101: color_data = 12'b111011101110;
20'b00100100110110101110: color_data = 12'b111011101110;
20'b00100100110110101111: color_data = 12'b111011101110;
20'b00100100110110110000: color_data = 12'b111011101110;
20'b00100100110110110001: color_data = 12'b111011101110;
20'b00100100110110110010: color_data = 12'b111011101110;
20'b00100100110110110100: color_data = 12'b111011101110;
20'b00100100110110110101: color_data = 12'b111011101110;
20'b00100100110110110110: color_data = 12'b111011101110;
20'b00100100110110110111: color_data = 12'b111011101110;
20'b00100100110110111000: color_data = 12'b111011101110;
20'b00100100110110111001: color_data = 12'b111011101110;
20'b00100100110110111010: color_data = 12'b111011101110;
20'b00100100110110111011: color_data = 12'b111011101110;
20'b00100100110110111100: color_data = 12'b111011101110;
20'b00100100110110111101: color_data = 12'b111011101110;
20'b00100100110110111111: color_data = 12'b111011101110;
20'b00100100110111000000: color_data = 12'b111011101110;
20'b00100100110111000001: color_data = 12'b111011101110;
20'b00100100110111000010: color_data = 12'b111011101110;
20'b00100100110111000011: color_data = 12'b111011101110;
20'b00100100110111000100: color_data = 12'b111011101110;
20'b00100100110111000101: color_data = 12'b111011101110;
20'b00100100110111000110: color_data = 12'b111011101110;
20'b00100100110111000111: color_data = 12'b111011101110;
20'b00100100110111001000: color_data = 12'b111011101110;
20'b00100100110111001010: color_data = 12'b111011101110;
20'b00100100110111001011: color_data = 12'b111011101110;
20'b00100100110111001100: color_data = 12'b111011101110;
20'b00100100110111001101: color_data = 12'b111011101110;
20'b00100100110111001110: color_data = 12'b111011101110;
20'b00100100110111001111: color_data = 12'b111011101110;
20'b00100100110111010000: color_data = 12'b111011101110;
20'b00100100110111010001: color_data = 12'b111011101110;
20'b00100100110111010010: color_data = 12'b111011101110;
20'b00100100110111010011: color_data = 12'b111011101110;
20'b00100101000010010110: color_data = 12'b111011101110;
20'b00100101000010010111: color_data = 12'b111011101110;
20'b00100101000010011000: color_data = 12'b111011101110;
20'b00100101000010011001: color_data = 12'b111011101110;
20'b00100101000010011010: color_data = 12'b111011101110;
20'b00100101000010011011: color_data = 12'b111011101110;
20'b00100101000010011100: color_data = 12'b111011101110;
20'b00100101000010011101: color_data = 12'b111011101110;
20'b00100101000010011110: color_data = 12'b111011101110;
20'b00100101000010011111: color_data = 12'b111011101110;
20'b00100101000010100001: color_data = 12'b111011101110;
20'b00100101000010100010: color_data = 12'b111011101110;
20'b00100101000010100011: color_data = 12'b111011101110;
20'b00100101000010100100: color_data = 12'b111011101110;
20'b00100101000010100101: color_data = 12'b111011101110;
20'b00100101000010100110: color_data = 12'b111011101110;
20'b00100101000010100111: color_data = 12'b111011101110;
20'b00100101000010101000: color_data = 12'b111011101110;
20'b00100101000010101001: color_data = 12'b111011101110;
20'b00100101000010101010: color_data = 12'b111011101110;
20'b00100101000011101110: color_data = 12'b111011101110;
20'b00100101000011101111: color_data = 12'b111011101110;
20'b00100101000011110000: color_data = 12'b111011101110;
20'b00100101000011110001: color_data = 12'b111011101110;
20'b00100101000011110010: color_data = 12'b111011101110;
20'b00100101000011110011: color_data = 12'b111011101110;
20'b00100101000011110100: color_data = 12'b111011101110;
20'b00100101000011110101: color_data = 12'b111011101110;
20'b00100101000011110110: color_data = 12'b111011101110;
20'b00100101000011110111: color_data = 12'b111011101110;
20'b00100101000011111001: color_data = 12'b111011101110;
20'b00100101000011111010: color_data = 12'b111011101110;
20'b00100101000011111011: color_data = 12'b111011101110;
20'b00100101000011111100: color_data = 12'b111011101110;
20'b00100101000011111101: color_data = 12'b111011101110;
20'b00100101000011111110: color_data = 12'b111011101110;
20'b00100101000011111111: color_data = 12'b111011101110;
20'b00100101000100000000: color_data = 12'b111011101110;
20'b00100101000100000001: color_data = 12'b111011101110;
20'b00100101000100000010: color_data = 12'b111011101110;
20'b00100101000100100101: color_data = 12'b111011101110;
20'b00100101000100100110: color_data = 12'b111011101110;
20'b00100101000100100111: color_data = 12'b111011101110;
20'b00100101000100101000: color_data = 12'b111011101110;
20'b00100101000100101001: color_data = 12'b111011101110;
20'b00100101000100101010: color_data = 12'b111011101110;
20'b00100101000100101011: color_data = 12'b111011101110;
20'b00100101000100101100: color_data = 12'b111011101110;
20'b00100101000100101101: color_data = 12'b111011101110;
20'b00100101000100101110: color_data = 12'b111011101110;
20'b00100101000100110000: color_data = 12'b111011101110;
20'b00100101000100110001: color_data = 12'b111011101110;
20'b00100101000100110010: color_data = 12'b111011101110;
20'b00100101000100110011: color_data = 12'b111011101110;
20'b00100101000100110100: color_data = 12'b111011101110;
20'b00100101000100110101: color_data = 12'b111011101110;
20'b00100101000100110110: color_data = 12'b111011101110;
20'b00100101000100110111: color_data = 12'b111011101110;
20'b00100101000100111000: color_data = 12'b111011101110;
20'b00100101000100111001: color_data = 12'b111011101110;
20'b00100101000101000110: color_data = 12'b111011101110;
20'b00100101000101000111: color_data = 12'b111011101110;
20'b00100101000101001000: color_data = 12'b111011101110;
20'b00100101000101001001: color_data = 12'b111011101110;
20'b00100101000101001010: color_data = 12'b111011101110;
20'b00100101000101001011: color_data = 12'b111011101110;
20'b00100101000101001100: color_data = 12'b111011101110;
20'b00100101000101001101: color_data = 12'b111011101110;
20'b00100101000101001110: color_data = 12'b111011101110;
20'b00100101000101001111: color_data = 12'b111011101110;
20'b00100101000101010001: color_data = 12'b111011101110;
20'b00100101000101010010: color_data = 12'b111011101110;
20'b00100101000101010011: color_data = 12'b111011101110;
20'b00100101000101010100: color_data = 12'b111011101110;
20'b00100101000101010101: color_data = 12'b111011101110;
20'b00100101000101010110: color_data = 12'b111011101110;
20'b00100101000101010111: color_data = 12'b111011101110;
20'b00100101000101011000: color_data = 12'b111011101110;
20'b00100101000101011001: color_data = 12'b111011101110;
20'b00100101000101011010: color_data = 12'b111011101110;
20'b00100101000101100111: color_data = 12'b111011101110;
20'b00100101000101101000: color_data = 12'b111011101110;
20'b00100101000101101001: color_data = 12'b111011101110;
20'b00100101000101101010: color_data = 12'b111011101110;
20'b00100101000101101011: color_data = 12'b111011101110;
20'b00100101000101101100: color_data = 12'b111011101110;
20'b00100101000101101101: color_data = 12'b111011101110;
20'b00100101000101101110: color_data = 12'b111011101110;
20'b00100101000101101111: color_data = 12'b111011101110;
20'b00100101000101110000: color_data = 12'b111011101110;
20'b00100101000101111101: color_data = 12'b111011101110;
20'b00100101000101111110: color_data = 12'b111011101110;
20'b00100101000101111111: color_data = 12'b111011101110;
20'b00100101000110000000: color_data = 12'b111011101110;
20'b00100101000110000001: color_data = 12'b111011101110;
20'b00100101000110000010: color_data = 12'b111011101110;
20'b00100101000110000011: color_data = 12'b111011101110;
20'b00100101000110000100: color_data = 12'b111011101110;
20'b00100101000110000101: color_data = 12'b111011101110;
20'b00100101000110000110: color_data = 12'b111011101110;
20'b00100101000110001000: color_data = 12'b111011101110;
20'b00100101000110001001: color_data = 12'b111011101110;
20'b00100101000110001010: color_data = 12'b111011101110;
20'b00100101000110001011: color_data = 12'b111011101110;
20'b00100101000110001100: color_data = 12'b111011101110;
20'b00100101000110001101: color_data = 12'b111011101110;
20'b00100101000110001110: color_data = 12'b111011101110;
20'b00100101000110001111: color_data = 12'b111011101110;
20'b00100101000110010000: color_data = 12'b111011101110;
20'b00100101000110010001: color_data = 12'b111011101110;
20'b00100101000110011110: color_data = 12'b111011101110;
20'b00100101000110011111: color_data = 12'b111011101110;
20'b00100101000110100000: color_data = 12'b111011101110;
20'b00100101000110100001: color_data = 12'b111011101110;
20'b00100101000110100010: color_data = 12'b111011101110;
20'b00100101000110100011: color_data = 12'b111011101110;
20'b00100101000110100100: color_data = 12'b111011101110;
20'b00100101000110100101: color_data = 12'b111011101110;
20'b00100101000110100110: color_data = 12'b111011101110;
20'b00100101000110100111: color_data = 12'b111011101110;
20'b00100101000110101001: color_data = 12'b111011101110;
20'b00100101000110101010: color_data = 12'b111011101110;
20'b00100101000110101011: color_data = 12'b111011101110;
20'b00100101000110101100: color_data = 12'b111011101110;
20'b00100101000110101101: color_data = 12'b111011101110;
20'b00100101000110101110: color_data = 12'b111011101110;
20'b00100101000110101111: color_data = 12'b111011101110;
20'b00100101000110110000: color_data = 12'b111011101110;
20'b00100101000110110001: color_data = 12'b111011101110;
20'b00100101000110110010: color_data = 12'b111011101110;
20'b00100101000110110100: color_data = 12'b111011101110;
20'b00100101000110110101: color_data = 12'b111011101110;
20'b00100101000110110110: color_data = 12'b111011101110;
20'b00100101000110110111: color_data = 12'b111011101110;
20'b00100101000110111000: color_data = 12'b111011101110;
20'b00100101000110111001: color_data = 12'b111011101110;
20'b00100101000110111010: color_data = 12'b111011101110;
20'b00100101000110111011: color_data = 12'b111011101110;
20'b00100101000110111100: color_data = 12'b111011101110;
20'b00100101000110111101: color_data = 12'b111011101110;
20'b00100101000110111111: color_data = 12'b111011101110;
20'b00100101000111000000: color_data = 12'b111011101110;
20'b00100101000111000001: color_data = 12'b111011101110;
20'b00100101000111000010: color_data = 12'b111011101110;
20'b00100101000111000011: color_data = 12'b111011101110;
20'b00100101000111000100: color_data = 12'b111011101110;
20'b00100101000111000101: color_data = 12'b111011101110;
20'b00100101000111000110: color_data = 12'b111011101110;
20'b00100101000111000111: color_data = 12'b111011101110;
20'b00100101000111001000: color_data = 12'b111011101110;
20'b00100101000111001010: color_data = 12'b111011101110;
20'b00100101000111001011: color_data = 12'b111011101110;
20'b00100101000111001100: color_data = 12'b111011101110;
20'b00100101000111001101: color_data = 12'b111011101110;
20'b00100101000111001110: color_data = 12'b111011101110;
20'b00100101000111001111: color_data = 12'b111011101110;
20'b00100101000111010000: color_data = 12'b111011101110;
20'b00100101000111010001: color_data = 12'b111011101110;
20'b00100101000111010010: color_data = 12'b111011101110;
20'b00100101000111010011: color_data = 12'b111011101110;
20'b00100101010010010110: color_data = 12'b111011101110;
20'b00100101010010010111: color_data = 12'b111011101110;
20'b00100101010010011000: color_data = 12'b111011101110;
20'b00100101010010011001: color_data = 12'b111011101110;
20'b00100101010010011010: color_data = 12'b111011101110;
20'b00100101010010011011: color_data = 12'b111011101110;
20'b00100101010010011100: color_data = 12'b111011101110;
20'b00100101010010011101: color_data = 12'b111011101110;
20'b00100101010010011110: color_data = 12'b111011101110;
20'b00100101010010011111: color_data = 12'b111011101110;
20'b00100101010010100001: color_data = 12'b111011101110;
20'b00100101010010100010: color_data = 12'b111011101110;
20'b00100101010010100011: color_data = 12'b111011101110;
20'b00100101010010100100: color_data = 12'b111011101110;
20'b00100101010010100101: color_data = 12'b111011101110;
20'b00100101010010100110: color_data = 12'b111011101110;
20'b00100101010010100111: color_data = 12'b111011101110;
20'b00100101010010101000: color_data = 12'b111011101110;
20'b00100101010010101001: color_data = 12'b111011101110;
20'b00100101010010101010: color_data = 12'b111011101110;
20'b00100101010011101110: color_data = 12'b111011101110;
20'b00100101010011101111: color_data = 12'b111011101110;
20'b00100101010011110000: color_data = 12'b111011101110;
20'b00100101010011110001: color_data = 12'b111011101110;
20'b00100101010011110010: color_data = 12'b111011101110;
20'b00100101010011110011: color_data = 12'b111011101110;
20'b00100101010011110100: color_data = 12'b111011101110;
20'b00100101010011110101: color_data = 12'b111011101110;
20'b00100101010011110110: color_data = 12'b111011101110;
20'b00100101010011110111: color_data = 12'b111011101110;
20'b00100101010011111001: color_data = 12'b111011101110;
20'b00100101010011111010: color_data = 12'b111011101110;
20'b00100101010011111011: color_data = 12'b111011101110;
20'b00100101010011111100: color_data = 12'b111011101110;
20'b00100101010011111101: color_data = 12'b111011101110;
20'b00100101010011111110: color_data = 12'b111011101110;
20'b00100101010011111111: color_data = 12'b111011101110;
20'b00100101010100000000: color_data = 12'b111011101110;
20'b00100101010100000001: color_data = 12'b111011101110;
20'b00100101010100000010: color_data = 12'b111011101110;
20'b00100101010100100101: color_data = 12'b111011101110;
20'b00100101010100100110: color_data = 12'b111011101110;
20'b00100101010100100111: color_data = 12'b111011101110;
20'b00100101010100101000: color_data = 12'b111011101110;
20'b00100101010100101001: color_data = 12'b111011101110;
20'b00100101010100101010: color_data = 12'b111011101110;
20'b00100101010100101011: color_data = 12'b111011101110;
20'b00100101010100101100: color_data = 12'b111011101110;
20'b00100101010100101101: color_data = 12'b111011101110;
20'b00100101010100101110: color_data = 12'b111011101110;
20'b00100101010100110000: color_data = 12'b111011101110;
20'b00100101010100110001: color_data = 12'b111011101110;
20'b00100101010100110010: color_data = 12'b111011101110;
20'b00100101010100110011: color_data = 12'b111011101110;
20'b00100101010100110100: color_data = 12'b111011101110;
20'b00100101010100110101: color_data = 12'b111011101110;
20'b00100101010100110110: color_data = 12'b111011101110;
20'b00100101010100110111: color_data = 12'b111011101110;
20'b00100101010100111000: color_data = 12'b111011101110;
20'b00100101010100111001: color_data = 12'b111011101110;
20'b00100101010101000110: color_data = 12'b111011101110;
20'b00100101010101000111: color_data = 12'b111011101110;
20'b00100101010101001000: color_data = 12'b111011101110;
20'b00100101010101001001: color_data = 12'b111011101110;
20'b00100101010101001010: color_data = 12'b111011101110;
20'b00100101010101001011: color_data = 12'b111011101110;
20'b00100101010101001100: color_data = 12'b111011101110;
20'b00100101010101001101: color_data = 12'b111011101110;
20'b00100101010101001110: color_data = 12'b111011101110;
20'b00100101010101001111: color_data = 12'b111011101110;
20'b00100101010101010001: color_data = 12'b111011101110;
20'b00100101010101010010: color_data = 12'b111011101110;
20'b00100101010101010011: color_data = 12'b111011101110;
20'b00100101010101010100: color_data = 12'b111011101110;
20'b00100101010101010101: color_data = 12'b111011101110;
20'b00100101010101010110: color_data = 12'b111011101110;
20'b00100101010101010111: color_data = 12'b111011101110;
20'b00100101010101011000: color_data = 12'b111011101110;
20'b00100101010101011001: color_data = 12'b111011101110;
20'b00100101010101011010: color_data = 12'b111011101110;
20'b00100101010101100111: color_data = 12'b111011101110;
20'b00100101010101101000: color_data = 12'b111011101110;
20'b00100101010101101001: color_data = 12'b111011101110;
20'b00100101010101101010: color_data = 12'b111011101110;
20'b00100101010101101011: color_data = 12'b111011101110;
20'b00100101010101101100: color_data = 12'b111011101110;
20'b00100101010101101101: color_data = 12'b111011101110;
20'b00100101010101101110: color_data = 12'b111011101110;
20'b00100101010101101111: color_data = 12'b111011101110;
20'b00100101010101110000: color_data = 12'b111011101110;
20'b00100101010101111101: color_data = 12'b111011101110;
20'b00100101010101111110: color_data = 12'b111011101110;
20'b00100101010101111111: color_data = 12'b111011101110;
20'b00100101010110000000: color_data = 12'b111011101110;
20'b00100101010110000001: color_data = 12'b111011101110;
20'b00100101010110000010: color_data = 12'b111011101110;
20'b00100101010110000011: color_data = 12'b111011101110;
20'b00100101010110000100: color_data = 12'b111011101110;
20'b00100101010110000101: color_data = 12'b111011101110;
20'b00100101010110000110: color_data = 12'b111011101110;
20'b00100101010110001000: color_data = 12'b111011101110;
20'b00100101010110001001: color_data = 12'b111011101110;
20'b00100101010110001010: color_data = 12'b111011101110;
20'b00100101010110001011: color_data = 12'b111011101110;
20'b00100101010110001100: color_data = 12'b111011101110;
20'b00100101010110001101: color_data = 12'b111011101110;
20'b00100101010110001110: color_data = 12'b111011101110;
20'b00100101010110001111: color_data = 12'b111011101110;
20'b00100101010110010000: color_data = 12'b111011101110;
20'b00100101010110010001: color_data = 12'b111011101110;
20'b00100101010110011110: color_data = 12'b111011101110;
20'b00100101010110011111: color_data = 12'b111011101110;
20'b00100101010110100000: color_data = 12'b111011101110;
20'b00100101010110100001: color_data = 12'b111011101110;
20'b00100101010110100010: color_data = 12'b111011101110;
20'b00100101010110100011: color_data = 12'b111011101110;
20'b00100101010110100100: color_data = 12'b111011101110;
20'b00100101010110100101: color_data = 12'b111011101110;
20'b00100101010110100110: color_data = 12'b111011101110;
20'b00100101010110100111: color_data = 12'b111011101110;
20'b00100101010110101001: color_data = 12'b111011101110;
20'b00100101010110101010: color_data = 12'b111011101110;
20'b00100101010110101011: color_data = 12'b111011101110;
20'b00100101010110101100: color_data = 12'b111011101110;
20'b00100101010110101101: color_data = 12'b111011101110;
20'b00100101010110101110: color_data = 12'b111011101110;
20'b00100101010110101111: color_data = 12'b111011101110;
20'b00100101010110110000: color_data = 12'b111011101110;
20'b00100101010110110001: color_data = 12'b111011101110;
20'b00100101010110110010: color_data = 12'b111011101110;
20'b00100101010110110100: color_data = 12'b111011101110;
20'b00100101010110110101: color_data = 12'b111011101110;
20'b00100101010110110110: color_data = 12'b111011101110;
20'b00100101010110110111: color_data = 12'b111011101110;
20'b00100101010110111000: color_data = 12'b111011101110;
20'b00100101010110111001: color_data = 12'b111011101110;
20'b00100101010110111010: color_data = 12'b111011101110;
20'b00100101010110111011: color_data = 12'b111011101110;
20'b00100101010110111100: color_data = 12'b111011101110;
20'b00100101010110111101: color_data = 12'b111011101110;
20'b00100101010110111111: color_data = 12'b111011101110;
20'b00100101010111000000: color_data = 12'b111011101110;
20'b00100101010111000001: color_data = 12'b111011101110;
20'b00100101010111000010: color_data = 12'b111011101110;
20'b00100101010111000011: color_data = 12'b111011101110;
20'b00100101010111000100: color_data = 12'b111011101110;
20'b00100101010111000101: color_data = 12'b111011101110;
20'b00100101010111000110: color_data = 12'b111011101110;
20'b00100101010111000111: color_data = 12'b111011101110;
20'b00100101010111001000: color_data = 12'b111011101110;
20'b00100101010111001010: color_data = 12'b111011101110;
20'b00100101010111001011: color_data = 12'b111011101110;
20'b00100101010111001100: color_data = 12'b111011101110;
20'b00100101010111001101: color_data = 12'b111011101110;
20'b00100101010111001110: color_data = 12'b111011101110;
20'b00100101010111001111: color_data = 12'b111011101110;
20'b00100101010111010000: color_data = 12'b111011101110;
20'b00100101010111010001: color_data = 12'b111011101110;
20'b00100101010111010010: color_data = 12'b111011101110;
20'b00100101010111010011: color_data = 12'b111011101110;
20'b00100101100010010110: color_data = 12'b111011101110;
20'b00100101100010010111: color_data = 12'b111011101110;
20'b00100101100010011000: color_data = 12'b111011101110;
20'b00100101100010011001: color_data = 12'b111011101110;
20'b00100101100010011010: color_data = 12'b111011101110;
20'b00100101100010011011: color_data = 12'b111011101110;
20'b00100101100010011100: color_data = 12'b111011101110;
20'b00100101100010011101: color_data = 12'b111011101110;
20'b00100101100010011110: color_data = 12'b111011101110;
20'b00100101100010011111: color_data = 12'b111011101110;
20'b00100101100010100001: color_data = 12'b111011101110;
20'b00100101100010100010: color_data = 12'b111011101110;
20'b00100101100010100011: color_data = 12'b111011101110;
20'b00100101100010100100: color_data = 12'b111011101110;
20'b00100101100010100101: color_data = 12'b111011101110;
20'b00100101100010100110: color_data = 12'b111011101110;
20'b00100101100010100111: color_data = 12'b111011101110;
20'b00100101100010101000: color_data = 12'b111011101110;
20'b00100101100010101001: color_data = 12'b111011101110;
20'b00100101100010101010: color_data = 12'b111011101110;
20'b00100101100011101110: color_data = 12'b111011101110;
20'b00100101100011101111: color_data = 12'b111011101110;
20'b00100101100011110000: color_data = 12'b111011101110;
20'b00100101100011110001: color_data = 12'b111011101110;
20'b00100101100011110010: color_data = 12'b111011101110;
20'b00100101100011110011: color_data = 12'b111011101110;
20'b00100101100011110100: color_data = 12'b111011101110;
20'b00100101100011110101: color_data = 12'b111011101110;
20'b00100101100011110110: color_data = 12'b111011101110;
20'b00100101100011110111: color_data = 12'b111011101110;
20'b00100101100011111001: color_data = 12'b111011101110;
20'b00100101100011111010: color_data = 12'b111011101110;
20'b00100101100011111011: color_data = 12'b111011101110;
20'b00100101100011111100: color_data = 12'b111011101110;
20'b00100101100011111101: color_data = 12'b111011101110;
20'b00100101100011111110: color_data = 12'b111011101110;
20'b00100101100011111111: color_data = 12'b111011101110;
20'b00100101100100000000: color_data = 12'b111011101110;
20'b00100101100100000001: color_data = 12'b111011101110;
20'b00100101100100000010: color_data = 12'b111011101110;
20'b00100101100100100101: color_data = 12'b111011101110;
20'b00100101100100100110: color_data = 12'b111011101110;
20'b00100101100100100111: color_data = 12'b111011101110;
20'b00100101100100101000: color_data = 12'b111011101110;
20'b00100101100100101001: color_data = 12'b111011101110;
20'b00100101100100101010: color_data = 12'b111011101110;
20'b00100101100100101011: color_data = 12'b111011101110;
20'b00100101100100101100: color_data = 12'b111011101110;
20'b00100101100100101101: color_data = 12'b111011101110;
20'b00100101100100101110: color_data = 12'b111011101110;
20'b00100101100100110000: color_data = 12'b111011101110;
20'b00100101100100110001: color_data = 12'b111011101110;
20'b00100101100100110010: color_data = 12'b111011101110;
20'b00100101100100110011: color_data = 12'b111011101110;
20'b00100101100100110100: color_data = 12'b111011101110;
20'b00100101100100110101: color_data = 12'b111011101110;
20'b00100101100100110110: color_data = 12'b111011101110;
20'b00100101100100110111: color_data = 12'b111011101110;
20'b00100101100100111000: color_data = 12'b111011101110;
20'b00100101100100111001: color_data = 12'b111011101110;
20'b00100101100101000110: color_data = 12'b111011101110;
20'b00100101100101000111: color_data = 12'b111011101110;
20'b00100101100101001000: color_data = 12'b111011101110;
20'b00100101100101001001: color_data = 12'b111011101110;
20'b00100101100101001010: color_data = 12'b111011101110;
20'b00100101100101001011: color_data = 12'b111011101110;
20'b00100101100101001100: color_data = 12'b111011101110;
20'b00100101100101001101: color_data = 12'b111011101110;
20'b00100101100101001110: color_data = 12'b111011101110;
20'b00100101100101001111: color_data = 12'b111011101110;
20'b00100101100101010001: color_data = 12'b111011101110;
20'b00100101100101010010: color_data = 12'b111011101110;
20'b00100101100101010011: color_data = 12'b111011101110;
20'b00100101100101010100: color_data = 12'b111011101110;
20'b00100101100101010101: color_data = 12'b111011101110;
20'b00100101100101010110: color_data = 12'b111011101110;
20'b00100101100101010111: color_data = 12'b111011101110;
20'b00100101100101011000: color_data = 12'b111011101110;
20'b00100101100101011001: color_data = 12'b111011101110;
20'b00100101100101011010: color_data = 12'b111011101110;
20'b00100101100101100111: color_data = 12'b111011101110;
20'b00100101100101101000: color_data = 12'b111011101110;
20'b00100101100101101001: color_data = 12'b111011101110;
20'b00100101100101101010: color_data = 12'b111011101110;
20'b00100101100101101011: color_data = 12'b111011101110;
20'b00100101100101101100: color_data = 12'b111011101110;
20'b00100101100101101101: color_data = 12'b111011101110;
20'b00100101100101101110: color_data = 12'b111011101110;
20'b00100101100101101111: color_data = 12'b111011101110;
20'b00100101100101110000: color_data = 12'b111011101110;
20'b00100101100101111101: color_data = 12'b111011101110;
20'b00100101100101111110: color_data = 12'b111011101110;
20'b00100101100101111111: color_data = 12'b111011101110;
20'b00100101100110000000: color_data = 12'b111011101110;
20'b00100101100110000001: color_data = 12'b111011101110;
20'b00100101100110000010: color_data = 12'b111011101110;
20'b00100101100110000011: color_data = 12'b111011101110;
20'b00100101100110000100: color_data = 12'b111011101110;
20'b00100101100110000101: color_data = 12'b111011101110;
20'b00100101100110000110: color_data = 12'b111011101110;
20'b00100101100110001000: color_data = 12'b111011101110;
20'b00100101100110001001: color_data = 12'b111011101110;
20'b00100101100110001010: color_data = 12'b111011101110;
20'b00100101100110001011: color_data = 12'b111011101110;
20'b00100101100110001100: color_data = 12'b111011101110;
20'b00100101100110001101: color_data = 12'b111011101110;
20'b00100101100110001110: color_data = 12'b111011101110;
20'b00100101100110001111: color_data = 12'b111011101110;
20'b00100101100110010000: color_data = 12'b111011101110;
20'b00100101100110010001: color_data = 12'b111011101110;
20'b00100101100110011110: color_data = 12'b111011101110;
20'b00100101100110011111: color_data = 12'b111011101110;
20'b00100101100110100000: color_data = 12'b111011101110;
20'b00100101100110100001: color_data = 12'b111011101110;
20'b00100101100110100010: color_data = 12'b111011101110;
20'b00100101100110100011: color_data = 12'b111011101110;
20'b00100101100110100100: color_data = 12'b111011101110;
20'b00100101100110100101: color_data = 12'b111011101110;
20'b00100101100110100110: color_data = 12'b111011101110;
20'b00100101100110100111: color_data = 12'b111011101110;
20'b00100101100110101001: color_data = 12'b111011101110;
20'b00100101100110101010: color_data = 12'b111011101110;
20'b00100101100110101011: color_data = 12'b111011101110;
20'b00100101100110101100: color_data = 12'b111011101110;
20'b00100101100110101101: color_data = 12'b111011101110;
20'b00100101100110101110: color_data = 12'b111011101110;
20'b00100101100110101111: color_data = 12'b111011101110;
20'b00100101100110110000: color_data = 12'b111011101110;
20'b00100101100110110001: color_data = 12'b111011101110;
20'b00100101100110110010: color_data = 12'b111011101110;
20'b00100101100110110100: color_data = 12'b111011101110;
20'b00100101100110110101: color_data = 12'b111011101110;
20'b00100101100110110110: color_data = 12'b111011101110;
20'b00100101100110110111: color_data = 12'b111011101110;
20'b00100101100110111000: color_data = 12'b111011101110;
20'b00100101100110111001: color_data = 12'b111011101110;
20'b00100101100110111010: color_data = 12'b111011101110;
20'b00100101100110111011: color_data = 12'b111011101110;
20'b00100101100110111100: color_data = 12'b111011101110;
20'b00100101100110111101: color_data = 12'b111011101110;
20'b00100101100110111111: color_data = 12'b111011101110;
20'b00100101100111000000: color_data = 12'b111011101110;
20'b00100101100111000001: color_data = 12'b111011101110;
20'b00100101100111000010: color_data = 12'b111011101110;
20'b00100101100111000011: color_data = 12'b111011101110;
20'b00100101100111000100: color_data = 12'b111011101110;
20'b00100101100111000101: color_data = 12'b111011101110;
20'b00100101100111000110: color_data = 12'b111011101110;
20'b00100101100111000111: color_data = 12'b111011101110;
20'b00100101100111001000: color_data = 12'b111011101110;
20'b00100101100111001010: color_data = 12'b111011101110;
20'b00100101100111001011: color_data = 12'b111011101110;
20'b00100101100111001100: color_data = 12'b111011101110;
20'b00100101100111001101: color_data = 12'b111011101110;
20'b00100101100111001110: color_data = 12'b111011101110;
20'b00100101100111001111: color_data = 12'b111011101110;
20'b00100101100111010000: color_data = 12'b111011101110;
20'b00100101100111010001: color_data = 12'b111011101110;
20'b00100101100111010010: color_data = 12'b111011101110;
20'b00100101100111010011: color_data = 12'b111011101110;
20'b00100101110010010110: color_data = 12'b111011101110;
20'b00100101110010010111: color_data = 12'b111011101110;
20'b00100101110010011000: color_data = 12'b111011101110;
20'b00100101110010011001: color_data = 12'b111011101110;
20'b00100101110010011010: color_data = 12'b111011101110;
20'b00100101110010011011: color_data = 12'b111011101110;
20'b00100101110010011100: color_data = 12'b111011101110;
20'b00100101110010011101: color_data = 12'b111011101110;
20'b00100101110010011110: color_data = 12'b111011101110;
20'b00100101110010011111: color_data = 12'b111011101110;
20'b00100101110010100001: color_data = 12'b111011101110;
20'b00100101110010100010: color_data = 12'b111011101110;
20'b00100101110010100011: color_data = 12'b111011101110;
20'b00100101110010100100: color_data = 12'b111011101110;
20'b00100101110010100101: color_data = 12'b111011101110;
20'b00100101110010100110: color_data = 12'b111011101110;
20'b00100101110010100111: color_data = 12'b111011101110;
20'b00100101110010101000: color_data = 12'b111011101110;
20'b00100101110010101001: color_data = 12'b111011101110;
20'b00100101110010101010: color_data = 12'b111011101110;
20'b00100101110011101110: color_data = 12'b111011101110;
20'b00100101110011101111: color_data = 12'b111011101110;
20'b00100101110011110000: color_data = 12'b111011101110;
20'b00100101110011110001: color_data = 12'b111011101110;
20'b00100101110011110010: color_data = 12'b111011101110;
20'b00100101110011110011: color_data = 12'b111011101110;
20'b00100101110011110100: color_data = 12'b111011101110;
20'b00100101110011110101: color_data = 12'b111011101110;
20'b00100101110011110110: color_data = 12'b111011101110;
20'b00100101110011110111: color_data = 12'b111011101110;
20'b00100101110011111001: color_data = 12'b111011101110;
20'b00100101110011111010: color_data = 12'b111011101110;
20'b00100101110011111011: color_data = 12'b111011101110;
20'b00100101110011111100: color_data = 12'b111011101110;
20'b00100101110011111101: color_data = 12'b111011101110;
20'b00100101110011111110: color_data = 12'b111011101110;
20'b00100101110011111111: color_data = 12'b111011101110;
20'b00100101110100000000: color_data = 12'b111011101110;
20'b00100101110100000001: color_data = 12'b111011101110;
20'b00100101110100000010: color_data = 12'b111011101110;
20'b00100101110100100101: color_data = 12'b111011101110;
20'b00100101110100100110: color_data = 12'b111011101110;
20'b00100101110100100111: color_data = 12'b111011101110;
20'b00100101110100101000: color_data = 12'b111011101110;
20'b00100101110100101001: color_data = 12'b111011101110;
20'b00100101110100101010: color_data = 12'b111011101110;
20'b00100101110100101011: color_data = 12'b111011101110;
20'b00100101110100101100: color_data = 12'b111011101110;
20'b00100101110100101101: color_data = 12'b111011101110;
20'b00100101110100101110: color_data = 12'b111011101110;
20'b00100101110100110000: color_data = 12'b111011101110;
20'b00100101110100110001: color_data = 12'b111011101110;
20'b00100101110100110010: color_data = 12'b111011101110;
20'b00100101110100110011: color_data = 12'b111011101110;
20'b00100101110100110100: color_data = 12'b111011101110;
20'b00100101110100110101: color_data = 12'b111011101110;
20'b00100101110100110110: color_data = 12'b111011101110;
20'b00100101110100110111: color_data = 12'b111011101110;
20'b00100101110100111000: color_data = 12'b111011101110;
20'b00100101110100111001: color_data = 12'b111011101110;
20'b00100101110101000110: color_data = 12'b111011101110;
20'b00100101110101000111: color_data = 12'b111011101110;
20'b00100101110101001000: color_data = 12'b111011101110;
20'b00100101110101001001: color_data = 12'b111011101110;
20'b00100101110101001010: color_data = 12'b111011101110;
20'b00100101110101001011: color_data = 12'b111011101110;
20'b00100101110101001100: color_data = 12'b111011101110;
20'b00100101110101001101: color_data = 12'b111011101110;
20'b00100101110101001110: color_data = 12'b111011101110;
20'b00100101110101001111: color_data = 12'b111011101110;
20'b00100101110101010001: color_data = 12'b111011101110;
20'b00100101110101010010: color_data = 12'b111011101110;
20'b00100101110101010011: color_data = 12'b111011101110;
20'b00100101110101010100: color_data = 12'b111011101110;
20'b00100101110101010101: color_data = 12'b111011101110;
20'b00100101110101010110: color_data = 12'b111011101110;
20'b00100101110101010111: color_data = 12'b111011101110;
20'b00100101110101011000: color_data = 12'b111011101110;
20'b00100101110101011001: color_data = 12'b111011101110;
20'b00100101110101011010: color_data = 12'b111011101110;
20'b00100101110101100111: color_data = 12'b111011101110;
20'b00100101110101101000: color_data = 12'b111011101110;
20'b00100101110101101001: color_data = 12'b111011101110;
20'b00100101110101101010: color_data = 12'b111011101110;
20'b00100101110101101011: color_data = 12'b111011101110;
20'b00100101110101101100: color_data = 12'b111011101110;
20'b00100101110101101101: color_data = 12'b111011101110;
20'b00100101110101101110: color_data = 12'b111011101110;
20'b00100101110101101111: color_data = 12'b111011101110;
20'b00100101110101110000: color_data = 12'b111011101110;
20'b00100101110101111101: color_data = 12'b111011101110;
20'b00100101110101111110: color_data = 12'b111011101110;
20'b00100101110101111111: color_data = 12'b111011101110;
20'b00100101110110000000: color_data = 12'b111011101110;
20'b00100101110110000001: color_data = 12'b111011101110;
20'b00100101110110000010: color_data = 12'b111011101110;
20'b00100101110110000011: color_data = 12'b111011101110;
20'b00100101110110000100: color_data = 12'b111011101110;
20'b00100101110110000101: color_data = 12'b111011101110;
20'b00100101110110000110: color_data = 12'b111011101110;
20'b00100101110110001000: color_data = 12'b111011101110;
20'b00100101110110001001: color_data = 12'b111011101110;
20'b00100101110110001010: color_data = 12'b111011101110;
20'b00100101110110001011: color_data = 12'b111011101110;
20'b00100101110110001100: color_data = 12'b111011101110;
20'b00100101110110001101: color_data = 12'b111011101110;
20'b00100101110110001110: color_data = 12'b111011101110;
20'b00100101110110001111: color_data = 12'b111011101110;
20'b00100101110110010000: color_data = 12'b111011101110;
20'b00100101110110010001: color_data = 12'b111011101110;
20'b00100101110110011110: color_data = 12'b111011101110;
20'b00100101110110011111: color_data = 12'b111011101110;
20'b00100101110110100000: color_data = 12'b111011101110;
20'b00100101110110100001: color_data = 12'b111011101110;
20'b00100101110110100010: color_data = 12'b111011101110;
20'b00100101110110100011: color_data = 12'b111011101110;
20'b00100101110110100100: color_data = 12'b111011101110;
20'b00100101110110100101: color_data = 12'b111011101110;
20'b00100101110110100110: color_data = 12'b111011101110;
20'b00100101110110100111: color_data = 12'b111011101110;
20'b00100101110110101001: color_data = 12'b111011101110;
20'b00100101110110101010: color_data = 12'b111011101110;
20'b00100101110110101011: color_data = 12'b111011101110;
20'b00100101110110101100: color_data = 12'b111011101110;
20'b00100101110110101101: color_data = 12'b111011101110;
20'b00100101110110101110: color_data = 12'b111011101110;
20'b00100101110110101111: color_data = 12'b111011101110;
20'b00100101110110110000: color_data = 12'b111011101110;
20'b00100101110110110001: color_data = 12'b111011101110;
20'b00100101110110110010: color_data = 12'b111011101110;
20'b00100101110110110100: color_data = 12'b111011101110;
20'b00100101110110110101: color_data = 12'b111011101110;
20'b00100101110110110110: color_data = 12'b111011101110;
20'b00100101110110110111: color_data = 12'b111011101110;
20'b00100101110110111000: color_data = 12'b111011101110;
20'b00100101110110111001: color_data = 12'b111011101110;
20'b00100101110110111010: color_data = 12'b111011101110;
20'b00100101110110111011: color_data = 12'b111011101110;
20'b00100101110110111100: color_data = 12'b111011101110;
20'b00100101110110111101: color_data = 12'b111011101110;
20'b00100101110110111111: color_data = 12'b111011101110;
20'b00100101110111000000: color_data = 12'b111011101110;
20'b00100101110111000001: color_data = 12'b111011101110;
20'b00100101110111000010: color_data = 12'b111011101110;
20'b00100101110111000011: color_data = 12'b111011101110;
20'b00100101110111000100: color_data = 12'b111011101110;
20'b00100101110111000101: color_data = 12'b111011101110;
20'b00100101110111000110: color_data = 12'b111011101110;
20'b00100101110111000111: color_data = 12'b111011101110;
20'b00100101110111001000: color_data = 12'b111011101110;
20'b00100101110111001010: color_data = 12'b111011101110;
20'b00100101110111001011: color_data = 12'b111011101110;
20'b00100101110111001100: color_data = 12'b111011101110;
20'b00100101110111001101: color_data = 12'b111011101110;
20'b00100101110111001110: color_data = 12'b111011101110;
20'b00100101110111001111: color_data = 12'b111011101110;
20'b00100101110111010000: color_data = 12'b111011101110;
20'b00100101110111010001: color_data = 12'b111011101110;
20'b00100101110111010010: color_data = 12'b111011101110;
20'b00100101110111010011: color_data = 12'b111011101110;
20'b00100110000010010110: color_data = 12'b111011101110;
20'b00100110000010010111: color_data = 12'b111011101110;
20'b00100110000010011000: color_data = 12'b111011101110;
20'b00100110000010011001: color_data = 12'b111011101110;
20'b00100110000010011010: color_data = 12'b111011101110;
20'b00100110000010011011: color_data = 12'b111011101110;
20'b00100110000010011100: color_data = 12'b111011101110;
20'b00100110000010011101: color_data = 12'b111011101110;
20'b00100110000010011110: color_data = 12'b111011101110;
20'b00100110000010011111: color_data = 12'b111011101110;
20'b00100110000010100001: color_data = 12'b111011101110;
20'b00100110000010100010: color_data = 12'b111011101110;
20'b00100110000010100011: color_data = 12'b111011101110;
20'b00100110000010100100: color_data = 12'b111011101110;
20'b00100110000010100101: color_data = 12'b111011101110;
20'b00100110000010100110: color_data = 12'b111011101110;
20'b00100110000010100111: color_data = 12'b111011101110;
20'b00100110000010101000: color_data = 12'b111011101110;
20'b00100110000010101001: color_data = 12'b111011101110;
20'b00100110000010101010: color_data = 12'b111011101110;
20'b00100110000011101110: color_data = 12'b111011101110;
20'b00100110000011101111: color_data = 12'b111011101110;
20'b00100110000011110000: color_data = 12'b111011101110;
20'b00100110000011110001: color_data = 12'b111011101110;
20'b00100110000011110010: color_data = 12'b111011101110;
20'b00100110000011110011: color_data = 12'b111011101110;
20'b00100110000011110100: color_data = 12'b111011101110;
20'b00100110000011110101: color_data = 12'b111011101110;
20'b00100110000011110110: color_data = 12'b111011101110;
20'b00100110000011110111: color_data = 12'b111011101110;
20'b00100110000011111001: color_data = 12'b111011101110;
20'b00100110000011111010: color_data = 12'b111011101110;
20'b00100110000011111011: color_data = 12'b111011101110;
20'b00100110000011111100: color_data = 12'b111011101110;
20'b00100110000011111101: color_data = 12'b111011101110;
20'b00100110000011111110: color_data = 12'b111011101110;
20'b00100110000011111111: color_data = 12'b111011101110;
20'b00100110000100000000: color_data = 12'b111011101110;
20'b00100110000100000001: color_data = 12'b111011101110;
20'b00100110000100000010: color_data = 12'b111011101110;
20'b00100110000100100101: color_data = 12'b111011101110;
20'b00100110000100100110: color_data = 12'b111011101110;
20'b00100110000100100111: color_data = 12'b111011101110;
20'b00100110000100101000: color_data = 12'b111011101110;
20'b00100110000100101001: color_data = 12'b111011101110;
20'b00100110000100101010: color_data = 12'b111011101110;
20'b00100110000100101011: color_data = 12'b111011101110;
20'b00100110000100101100: color_data = 12'b111011101110;
20'b00100110000100101101: color_data = 12'b111011101110;
20'b00100110000100101110: color_data = 12'b111011101110;
20'b00100110000100110000: color_data = 12'b111011101110;
20'b00100110000100110001: color_data = 12'b111011101110;
20'b00100110000100110010: color_data = 12'b111011101110;
20'b00100110000100110011: color_data = 12'b111011101110;
20'b00100110000100110100: color_data = 12'b111011101110;
20'b00100110000100110101: color_data = 12'b111011101110;
20'b00100110000100110110: color_data = 12'b111011101110;
20'b00100110000100110111: color_data = 12'b111011101110;
20'b00100110000100111000: color_data = 12'b111011101110;
20'b00100110000100111001: color_data = 12'b111011101110;
20'b00100110000101000110: color_data = 12'b111011101110;
20'b00100110000101000111: color_data = 12'b111011101110;
20'b00100110000101001000: color_data = 12'b111011101110;
20'b00100110000101001001: color_data = 12'b111011101110;
20'b00100110000101001010: color_data = 12'b111011101110;
20'b00100110000101001011: color_data = 12'b111011101110;
20'b00100110000101001100: color_data = 12'b111011101110;
20'b00100110000101001101: color_data = 12'b111011101110;
20'b00100110000101001110: color_data = 12'b111011101110;
20'b00100110000101001111: color_data = 12'b111011101110;
20'b00100110000101010001: color_data = 12'b111011101110;
20'b00100110000101010010: color_data = 12'b111011101110;
20'b00100110000101010011: color_data = 12'b111011101110;
20'b00100110000101010100: color_data = 12'b111011101110;
20'b00100110000101010101: color_data = 12'b111011101110;
20'b00100110000101010110: color_data = 12'b111011101110;
20'b00100110000101010111: color_data = 12'b111011101110;
20'b00100110000101011000: color_data = 12'b111011101110;
20'b00100110000101011001: color_data = 12'b111011101110;
20'b00100110000101011010: color_data = 12'b111011101110;
20'b00100110000101100111: color_data = 12'b111011101110;
20'b00100110000101101000: color_data = 12'b111011101110;
20'b00100110000101101001: color_data = 12'b111011101110;
20'b00100110000101101010: color_data = 12'b111011101110;
20'b00100110000101101011: color_data = 12'b111011101110;
20'b00100110000101101100: color_data = 12'b111011101110;
20'b00100110000101101101: color_data = 12'b111011101110;
20'b00100110000101101110: color_data = 12'b111011101110;
20'b00100110000101101111: color_data = 12'b111011101110;
20'b00100110000101110000: color_data = 12'b111011101110;
20'b00100110000101111101: color_data = 12'b111011101110;
20'b00100110000101111110: color_data = 12'b111011101110;
20'b00100110000101111111: color_data = 12'b111011101110;
20'b00100110000110000000: color_data = 12'b111011101110;
20'b00100110000110000001: color_data = 12'b111011101110;
20'b00100110000110000010: color_data = 12'b111011101110;
20'b00100110000110000011: color_data = 12'b111011101110;
20'b00100110000110000100: color_data = 12'b111011101110;
20'b00100110000110000101: color_data = 12'b111011101110;
20'b00100110000110000110: color_data = 12'b111011101110;
20'b00100110000110001000: color_data = 12'b111011101110;
20'b00100110000110001001: color_data = 12'b111011101110;
20'b00100110000110001010: color_data = 12'b111011101110;
20'b00100110000110001011: color_data = 12'b111011101110;
20'b00100110000110001100: color_data = 12'b111011101110;
20'b00100110000110001101: color_data = 12'b111011101110;
20'b00100110000110001110: color_data = 12'b111011101110;
20'b00100110000110001111: color_data = 12'b111011101110;
20'b00100110000110010000: color_data = 12'b111011101110;
20'b00100110000110010001: color_data = 12'b111011101110;
20'b00100110000110011110: color_data = 12'b111011101110;
20'b00100110000110011111: color_data = 12'b111011101110;
20'b00100110000110100000: color_data = 12'b111011101110;
20'b00100110000110100001: color_data = 12'b111011101110;
20'b00100110000110100010: color_data = 12'b111011101110;
20'b00100110000110100011: color_data = 12'b111011101110;
20'b00100110000110100100: color_data = 12'b111011101110;
20'b00100110000110100101: color_data = 12'b111011101110;
20'b00100110000110100110: color_data = 12'b111011101110;
20'b00100110000110100111: color_data = 12'b111011101110;
20'b00100110000110101001: color_data = 12'b111011101110;
20'b00100110000110101010: color_data = 12'b111011101110;
20'b00100110000110101011: color_data = 12'b111011101110;
20'b00100110000110101100: color_data = 12'b111011101110;
20'b00100110000110101101: color_data = 12'b111011101110;
20'b00100110000110101110: color_data = 12'b111011101110;
20'b00100110000110101111: color_data = 12'b111011101110;
20'b00100110000110110000: color_data = 12'b111011101110;
20'b00100110000110110001: color_data = 12'b111011101110;
20'b00100110000110110010: color_data = 12'b111011101110;
20'b00100110000110110100: color_data = 12'b111011101110;
20'b00100110000110110101: color_data = 12'b111011101110;
20'b00100110000110110110: color_data = 12'b111011101110;
20'b00100110000110110111: color_data = 12'b111011101110;
20'b00100110000110111000: color_data = 12'b111011101110;
20'b00100110000110111001: color_data = 12'b111011101110;
20'b00100110000110111010: color_data = 12'b111011101110;
20'b00100110000110111011: color_data = 12'b111011101110;
20'b00100110000110111100: color_data = 12'b111011101110;
20'b00100110000110111101: color_data = 12'b111011101110;
20'b00100110000110111111: color_data = 12'b111011101110;
20'b00100110000111000000: color_data = 12'b111011101110;
20'b00100110000111000001: color_data = 12'b111011101110;
20'b00100110000111000010: color_data = 12'b111011101110;
20'b00100110000111000011: color_data = 12'b111011101110;
20'b00100110000111000100: color_data = 12'b111011101110;
20'b00100110000111000101: color_data = 12'b111011101110;
20'b00100110000111000110: color_data = 12'b111011101110;
20'b00100110000111000111: color_data = 12'b111011101110;
20'b00100110000111001000: color_data = 12'b111011101110;
20'b00100110000111001010: color_data = 12'b111011101110;
20'b00100110000111001011: color_data = 12'b111011101110;
20'b00100110000111001100: color_data = 12'b111011101110;
20'b00100110000111001101: color_data = 12'b111011101110;
20'b00100110000111001110: color_data = 12'b111011101110;
20'b00100110000111001111: color_data = 12'b111011101110;
20'b00100110000111010000: color_data = 12'b111011101110;
20'b00100110000111010001: color_data = 12'b111011101110;
20'b00100110000111010010: color_data = 12'b111011101110;
20'b00100110000111010011: color_data = 12'b111011101110;
20'b00100110010010010110: color_data = 12'b111011101110;
20'b00100110010010010111: color_data = 12'b111011101110;
20'b00100110010010011000: color_data = 12'b111011101110;
20'b00100110010010011001: color_data = 12'b111011101110;
20'b00100110010010011010: color_data = 12'b111011101110;
20'b00100110010010011011: color_data = 12'b111011101110;
20'b00100110010010011100: color_data = 12'b111011101110;
20'b00100110010010011101: color_data = 12'b111011101110;
20'b00100110010010011110: color_data = 12'b111011101110;
20'b00100110010010011111: color_data = 12'b111011101110;
20'b00100110010010100001: color_data = 12'b111011101110;
20'b00100110010010100010: color_data = 12'b111011101110;
20'b00100110010010100011: color_data = 12'b111011101110;
20'b00100110010010100100: color_data = 12'b111011101110;
20'b00100110010010100101: color_data = 12'b111011101110;
20'b00100110010010100110: color_data = 12'b111011101110;
20'b00100110010010100111: color_data = 12'b111011101110;
20'b00100110010010101000: color_data = 12'b111011101110;
20'b00100110010010101001: color_data = 12'b111011101110;
20'b00100110010010101010: color_data = 12'b111011101110;
20'b00100110010011101110: color_data = 12'b111011101110;
20'b00100110010011101111: color_data = 12'b111011101110;
20'b00100110010011110000: color_data = 12'b111011101110;
20'b00100110010011110001: color_data = 12'b111011101110;
20'b00100110010011110010: color_data = 12'b111011101110;
20'b00100110010011110011: color_data = 12'b111011101110;
20'b00100110010011110100: color_data = 12'b111011101110;
20'b00100110010011110101: color_data = 12'b111011101110;
20'b00100110010011110110: color_data = 12'b111011101110;
20'b00100110010011110111: color_data = 12'b111011101110;
20'b00100110010011111001: color_data = 12'b111011101110;
20'b00100110010011111010: color_data = 12'b111011101110;
20'b00100110010011111011: color_data = 12'b111011101110;
20'b00100110010011111100: color_data = 12'b111011101110;
20'b00100110010011111101: color_data = 12'b111011101110;
20'b00100110010011111110: color_data = 12'b111011101110;
20'b00100110010011111111: color_data = 12'b111011101110;
20'b00100110010100000000: color_data = 12'b111011101110;
20'b00100110010100000001: color_data = 12'b111011101110;
20'b00100110010100000010: color_data = 12'b111011101110;
20'b00100110010100100101: color_data = 12'b111011101110;
20'b00100110010100100110: color_data = 12'b111011101110;
20'b00100110010100100111: color_data = 12'b111011101110;
20'b00100110010100101000: color_data = 12'b111011101110;
20'b00100110010100101001: color_data = 12'b111011101110;
20'b00100110010100101010: color_data = 12'b111011101110;
20'b00100110010100101011: color_data = 12'b111011101110;
20'b00100110010100101100: color_data = 12'b111011101110;
20'b00100110010100101101: color_data = 12'b111011101110;
20'b00100110010100101110: color_data = 12'b111011101110;
20'b00100110010100110000: color_data = 12'b111011101110;
20'b00100110010100110001: color_data = 12'b111011101110;
20'b00100110010100110010: color_data = 12'b111011101110;
20'b00100110010100110011: color_data = 12'b111011101110;
20'b00100110010100110100: color_data = 12'b111011101110;
20'b00100110010100110101: color_data = 12'b111011101110;
20'b00100110010100110110: color_data = 12'b111011101110;
20'b00100110010100110111: color_data = 12'b111011101110;
20'b00100110010100111000: color_data = 12'b111011101110;
20'b00100110010100111001: color_data = 12'b111011101110;
20'b00100110010101000110: color_data = 12'b111011101110;
20'b00100110010101000111: color_data = 12'b111011101110;
20'b00100110010101001000: color_data = 12'b111011101110;
20'b00100110010101001001: color_data = 12'b111011101110;
20'b00100110010101001010: color_data = 12'b111011101110;
20'b00100110010101001011: color_data = 12'b111011101110;
20'b00100110010101001100: color_data = 12'b111011101110;
20'b00100110010101001101: color_data = 12'b111011101110;
20'b00100110010101001110: color_data = 12'b111011101110;
20'b00100110010101001111: color_data = 12'b111011101110;
20'b00100110010101010001: color_data = 12'b111011101110;
20'b00100110010101010010: color_data = 12'b111011101110;
20'b00100110010101010011: color_data = 12'b111011101110;
20'b00100110010101010100: color_data = 12'b111011101110;
20'b00100110010101010101: color_data = 12'b111011101110;
20'b00100110010101010110: color_data = 12'b111011101110;
20'b00100110010101010111: color_data = 12'b111011101110;
20'b00100110010101011000: color_data = 12'b111011101110;
20'b00100110010101011001: color_data = 12'b111011101110;
20'b00100110010101011010: color_data = 12'b111011101110;
20'b00100110010101100111: color_data = 12'b111011101110;
20'b00100110010101101000: color_data = 12'b111011101110;
20'b00100110010101101001: color_data = 12'b111011101110;
20'b00100110010101101010: color_data = 12'b111011101110;
20'b00100110010101101011: color_data = 12'b111011101110;
20'b00100110010101101100: color_data = 12'b111011101110;
20'b00100110010101101101: color_data = 12'b111011101110;
20'b00100110010101101110: color_data = 12'b111011101110;
20'b00100110010101101111: color_data = 12'b111011101110;
20'b00100110010101110000: color_data = 12'b111011101110;
20'b00100110010101111101: color_data = 12'b111011101110;
20'b00100110010101111110: color_data = 12'b111011101110;
20'b00100110010101111111: color_data = 12'b111011101110;
20'b00100110010110000000: color_data = 12'b111011101110;
20'b00100110010110000001: color_data = 12'b111011101110;
20'b00100110010110000010: color_data = 12'b111011101110;
20'b00100110010110000011: color_data = 12'b111011101110;
20'b00100110010110000100: color_data = 12'b111011101110;
20'b00100110010110000101: color_data = 12'b111011101110;
20'b00100110010110000110: color_data = 12'b111011101110;
20'b00100110010110001000: color_data = 12'b111011101110;
20'b00100110010110001001: color_data = 12'b111011101110;
20'b00100110010110001010: color_data = 12'b111011101110;
20'b00100110010110001011: color_data = 12'b111011101110;
20'b00100110010110001100: color_data = 12'b111011101110;
20'b00100110010110001101: color_data = 12'b111011101110;
20'b00100110010110001110: color_data = 12'b111011101110;
20'b00100110010110001111: color_data = 12'b111011101110;
20'b00100110010110010000: color_data = 12'b111011101110;
20'b00100110010110010001: color_data = 12'b111011101110;
20'b00100110010110011110: color_data = 12'b111011101110;
20'b00100110010110011111: color_data = 12'b111011101110;
20'b00100110010110100000: color_data = 12'b111011101110;
20'b00100110010110100001: color_data = 12'b111011101110;
20'b00100110010110100010: color_data = 12'b111011101110;
20'b00100110010110100011: color_data = 12'b111011101110;
20'b00100110010110100100: color_data = 12'b111011101110;
20'b00100110010110100101: color_data = 12'b111011101110;
20'b00100110010110100110: color_data = 12'b111011101110;
20'b00100110010110100111: color_data = 12'b111011101110;
20'b00100110010110101001: color_data = 12'b111011101110;
20'b00100110010110101010: color_data = 12'b111011101110;
20'b00100110010110101011: color_data = 12'b111011101110;
20'b00100110010110101100: color_data = 12'b111011101110;
20'b00100110010110101101: color_data = 12'b111011101110;
20'b00100110010110101110: color_data = 12'b111011101110;
20'b00100110010110101111: color_data = 12'b111011101110;
20'b00100110010110110000: color_data = 12'b111011101110;
20'b00100110010110110001: color_data = 12'b111011101110;
20'b00100110010110110010: color_data = 12'b111011101110;
20'b00100110010110110100: color_data = 12'b111011101110;
20'b00100110010110110101: color_data = 12'b111011101110;
20'b00100110010110110110: color_data = 12'b111011101110;
20'b00100110010110110111: color_data = 12'b111011101110;
20'b00100110010110111000: color_data = 12'b111011101110;
20'b00100110010110111001: color_data = 12'b111011101110;
20'b00100110010110111010: color_data = 12'b111011101110;
20'b00100110010110111011: color_data = 12'b111011101110;
20'b00100110010110111100: color_data = 12'b111011101110;
20'b00100110010110111101: color_data = 12'b111011101110;
20'b00100110010110111111: color_data = 12'b111011101110;
20'b00100110010111000000: color_data = 12'b111011101110;
20'b00100110010111000001: color_data = 12'b111011101110;
20'b00100110010111000010: color_data = 12'b111011101110;
20'b00100110010111000011: color_data = 12'b111011101110;
20'b00100110010111000100: color_data = 12'b111011101110;
20'b00100110010111000101: color_data = 12'b111011101110;
20'b00100110010111000110: color_data = 12'b111011101110;
20'b00100110010111000111: color_data = 12'b111011101110;
20'b00100110010111001000: color_data = 12'b111011101110;
20'b00100110010111001010: color_data = 12'b111011101110;
20'b00100110010111001011: color_data = 12'b111011101110;
20'b00100110010111001100: color_data = 12'b111011101110;
20'b00100110010111001101: color_data = 12'b111011101110;
20'b00100110010111001110: color_data = 12'b111011101110;
20'b00100110010111001111: color_data = 12'b111011101110;
20'b00100110010111010000: color_data = 12'b111011101110;
20'b00100110010111010001: color_data = 12'b111011101110;
20'b00100110010111010010: color_data = 12'b111011101110;
20'b00100110010111010011: color_data = 12'b111011101110;
20'b00100110100010010110: color_data = 12'b111011101110;
20'b00100110100010010111: color_data = 12'b111011101110;
20'b00100110100010011000: color_data = 12'b111011101110;
20'b00100110100010011001: color_data = 12'b111011101110;
20'b00100110100010011010: color_data = 12'b111011101110;
20'b00100110100010011011: color_data = 12'b111011101110;
20'b00100110100010011100: color_data = 12'b111011101110;
20'b00100110100010011101: color_data = 12'b111011101110;
20'b00100110100010011110: color_data = 12'b111011101110;
20'b00100110100010011111: color_data = 12'b111011101110;
20'b00100110100010100001: color_data = 12'b111011101110;
20'b00100110100010100010: color_data = 12'b111011101110;
20'b00100110100010100011: color_data = 12'b111011101110;
20'b00100110100010100100: color_data = 12'b111011101110;
20'b00100110100010100101: color_data = 12'b111011101110;
20'b00100110100010100110: color_data = 12'b111011101110;
20'b00100110100010100111: color_data = 12'b111011101110;
20'b00100110100010101000: color_data = 12'b111011101110;
20'b00100110100010101001: color_data = 12'b111011101110;
20'b00100110100010101010: color_data = 12'b111011101110;
20'b00100110100011101110: color_data = 12'b111011101110;
20'b00100110100011101111: color_data = 12'b111011101110;
20'b00100110100011110000: color_data = 12'b111011101110;
20'b00100110100011110001: color_data = 12'b111011101110;
20'b00100110100011110010: color_data = 12'b111011101110;
20'b00100110100011110011: color_data = 12'b111011101110;
20'b00100110100011110100: color_data = 12'b111011101110;
20'b00100110100011110101: color_data = 12'b111011101110;
20'b00100110100011110110: color_data = 12'b111011101110;
20'b00100110100011110111: color_data = 12'b111011101110;
20'b00100110100011111001: color_data = 12'b111011101110;
20'b00100110100011111010: color_data = 12'b111011101110;
20'b00100110100011111011: color_data = 12'b111011101110;
20'b00100110100011111100: color_data = 12'b111011101110;
20'b00100110100011111101: color_data = 12'b111011101110;
20'b00100110100011111110: color_data = 12'b111011101110;
20'b00100110100011111111: color_data = 12'b111011101110;
20'b00100110100100000000: color_data = 12'b111011101110;
20'b00100110100100000001: color_data = 12'b111011101110;
20'b00100110100100000010: color_data = 12'b111011101110;
20'b00100110100100100101: color_data = 12'b111011101110;
20'b00100110100100100110: color_data = 12'b111011101110;
20'b00100110100100100111: color_data = 12'b111011101110;
20'b00100110100100101000: color_data = 12'b111011101110;
20'b00100110100100101001: color_data = 12'b111011101110;
20'b00100110100100101010: color_data = 12'b111011101110;
20'b00100110100100101011: color_data = 12'b111011101110;
20'b00100110100100101100: color_data = 12'b111011101110;
20'b00100110100100101101: color_data = 12'b111011101110;
20'b00100110100100101110: color_data = 12'b111011101110;
20'b00100110100100110000: color_data = 12'b111011101110;
20'b00100110100100110001: color_data = 12'b111011101110;
20'b00100110100100110010: color_data = 12'b111011101110;
20'b00100110100100110011: color_data = 12'b111011101110;
20'b00100110100100110100: color_data = 12'b111011101110;
20'b00100110100100110101: color_data = 12'b111011101110;
20'b00100110100100110110: color_data = 12'b111011101110;
20'b00100110100100110111: color_data = 12'b111011101110;
20'b00100110100100111000: color_data = 12'b111011101110;
20'b00100110100100111001: color_data = 12'b111011101110;
20'b00100110100101000110: color_data = 12'b111011101110;
20'b00100110100101000111: color_data = 12'b111011101110;
20'b00100110100101001000: color_data = 12'b111011101110;
20'b00100110100101001001: color_data = 12'b111011101110;
20'b00100110100101001010: color_data = 12'b111011101110;
20'b00100110100101001011: color_data = 12'b111011101110;
20'b00100110100101001100: color_data = 12'b111011101110;
20'b00100110100101001101: color_data = 12'b111011101110;
20'b00100110100101001110: color_data = 12'b111011101110;
20'b00100110100101001111: color_data = 12'b111011101110;
20'b00100110100101010001: color_data = 12'b111011101110;
20'b00100110100101010010: color_data = 12'b111011101110;
20'b00100110100101010011: color_data = 12'b111011101110;
20'b00100110100101010100: color_data = 12'b111011101110;
20'b00100110100101010101: color_data = 12'b111011101110;
20'b00100110100101010110: color_data = 12'b111011101110;
20'b00100110100101010111: color_data = 12'b111011101110;
20'b00100110100101011000: color_data = 12'b111011101110;
20'b00100110100101011001: color_data = 12'b111011101110;
20'b00100110100101011010: color_data = 12'b111011101110;
20'b00100110100101100111: color_data = 12'b111011101110;
20'b00100110100101101000: color_data = 12'b111011101110;
20'b00100110100101101001: color_data = 12'b111011101110;
20'b00100110100101101010: color_data = 12'b111011101110;
20'b00100110100101101011: color_data = 12'b111011101110;
20'b00100110100101101100: color_data = 12'b111011101110;
20'b00100110100101101101: color_data = 12'b111011101110;
20'b00100110100101101110: color_data = 12'b111011101110;
20'b00100110100101101111: color_data = 12'b111011101110;
20'b00100110100101110000: color_data = 12'b111011101110;
20'b00100110100101111101: color_data = 12'b111011101110;
20'b00100110100101111110: color_data = 12'b111011101110;
20'b00100110100101111111: color_data = 12'b111011101110;
20'b00100110100110000000: color_data = 12'b111011101110;
20'b00100110100110000001: color_data = 12'b111011101110;
20'b00100110100110000010: color_data = 12'b111011101110;
20'b00100110100110000011: color_data = 12'b111011101110;
20'b00100110100110000100: color_data = 12'b111011101110;
20'b00100110100110000101: color_data = 12'b111011101110;
20'b00100110100110000110: color_data = 12'b111011101110;
20'b00100110100110001000: color_data = 12'b111011101110;
20'b00100110100110001001: color_data = 12'b111011101110;
20'b00100110100110001010: color_data = 12'b111011101110;
20'b00100110100110001011: color_data = 12'b111011101110;
20'b00100110100110001100: color_data = 12'b111011101110;
20'b00100110100110001101: color_data = 12'b111011101110;
20'b00100110100110001110: color_data = 12'b111011101110;
20'b00100110100110001111: color_data = 12'b111011101110;
20'b00100110100110010000: color_data = 12'b111011101110;
20'b00100110100110010001: color_data = 12'b111011101110;
20'b00100110100110011110: color_data = 12'b111011101110;
20'b00100110100110011111: color_data = 12'b111011101110;
20'b00100110100110100000: color_data = 12'b111011101110;
20'b00100110100110100001: color_data = 12'b111011101110;
20'b00100110100110100010: color_data = 12'b111011101110;
20'b00100110100110100011: color_data = 12'b111011101110;
20'b00100110100110100100: color_data = 12'b111011101110;
20'b00100110100110100101: color_data = 12'b111011101110;
20'b00100110100110100110: color_data = 12'b111011101110;
20'b00100110100110100111: color_data = 12'b111011101110;
20'b00100110100110101001: color_data = 12'b111011101110;
20'b00100110100110101010: color_data = 12'b111011101110;
20'b00100110100110101011: color_data = 12'b111011101110;
20'b00100110100110101100: color_data = 12'b111011101110;
20'b00100110100110101101: color_data = 12'b111011101110;
20'b00100110100110101110: color_data = 12'b111011101110;
20'b00100110100110101111: color_data = 12'b111011101110;
20'b00100110100110110000: color_data = 12'b111011101110;
20'b00100110100110110001: color_data = 12'b111011101110;
20'b00100110100110110010: color_data = 12'b111011101110;
20'b00100110100110110100: color_data = 12'b111011101110;
20'b00100110100110110101: color_data = 12'b111011101110;
20'b00100110100110110110: color_data = 12'b111011101110;
20'b00100110100110110111: color_data = 12'b111011101110;
20'b00100110100110111000: color_data = 12'b111011101110;
20'b00100110100110111001: color_data = 12'b111011101110;
20'b00100110100110111010: color_data = 12'b111011101110;
20'b00100110100110111011: color_data = 12'b111011101110;
20'b00100110100110111100: color_data = 12'b111011101110;
20'b00100110100110111101: color_data = 12'b111011101110;
20'b00100110100110111111: color_data = 12'b111011101110;
20'b00100110100111000000: color_data = 12'b111011101110;
20'b00100110100111000001: color_data = 12'b111011101110;
20'b00100110100111000010: color_data = 12'b111011101110;
20'b00100110100111000011: color_data = 12'b111011101110;
20'b00100110100111000100: color_data = 12'b111011101110;
20'b00100110100111000101: color_data = 12'b111011101110;
20'b00100110100111000110: color_data = 12'b111011101110;
20'b00100110100111000111: color_data = 12'b111011101110;
20'b00100110100111001000: color_data = 12'b111011101110;
20'b00100110100111001010: color_data = 12'b111011101110;
20'b00100110100111001011: color_data = 12'b111011101110;
20'b00100110100111001100: color_data = 12'b111011101110;
20'b00100110100111001101: color_data = 12'b111011101110;
20'b00100110100111001110: color_data = 12'b111011101110;
20'b00100110100111001111: color_data = 12'b111011101110;
20'b00100110100111010000: color_data = 12'b111011101110;
20'b00100110100111010001: color_data = 12'b111011101110;
20'b00100110100111010010: color_data = 12'b111011101110;
20'b00100110100111010011: color_data = 12'b111011101110;
20'b00100110110010010110: color_data = 12'b111011101110;
20'b00100110110010010111: color_data = 12'b111011101110;
20'b00100110110010011000: color_data = 12'b111011101110;
20'b00100110110010011001: color_data = 12'b111011101110;
20'b00100110110010011010: color_data = 12'b111011101110;
20'b00100110110010011011: color_data = 12'b111011101110;
20'b00100110110010011100: color_data = 12'b111011101110;
20'b00100110110010011101: color_data = 12'b111011101110;
20'b00100110110010011110: color_data = 12'b111011101110;
20'b00100110110010011111: color_data = 12'b111011101110;
20'b00100110110010100001: color_data = 12'b111011101110;
20'b00100110110010100010: color_data = 12'b111011101110;
20'b00100110110010100011: color_data = 12'b111011101110;
20'b00100110110010100100: color_data = 12'b111011101110;
20'b00100110110010100101: color_data = 12'b111011101110;
20'b00100110110010100110: color_data = 12'b111011101110;
20'b00100110110010100111: color_data = 12'b111011101110;
20'b00100110110010101000: color_data = 12'b111011101110;
20'b00100110110010101001: color_data = 12'b111011101110;
20'b00100110110010101010: color_data = 12'b111011101110;
20'b00100110110011000010: color_data = 12'b111011101110;
20'b00100110110011000011: color_data = 12'b111011101110;
20'b00100110110011000100: color_data = 12'b111011101110;
20'b00100110110011000101: color_data = 12'b111011101110;
20'b00100110110011000110: color_data = 12'b111011101110;
20'b00100110110011000111: color_data = 12'b111011101110;
20'b00100110110011001000: color_data = 12'b111011101110;
20'b00100110110011001001: color_data = 12'b111011101110;
20'b00100110110011001010: color_data = 12'b111011101110;
20'b00100110110011001011: color_data = 12'b111011101110;
20'b00100110110011001101: color_data = 12'b111011101110;
20'b00100110110011001110: color_data = 12'b111011101110;
20'b00100110110011001111: color_data = 12'b111011101110;
20'b00100110110011010000: color_data = 12'b111011101110;
20'b00100110110011010001: color_data = 12'b111011101110;
20'b00100110110011010010: color_data = 12'b111011101110;
20'b00100110110011010011: color_data = 12'b111011101110;
20'b00100110110011010100: color_data = 12'b111011101110;
20'b00100110110011010101: color_data = 12'b111011101110;
20'b00100110110011010110: color_data = 12'b111011101110;
20'b00100110110011011000: color_data = 12'b111011101110;
20'b00100110110011011001: color_data = 12'b111011101110;
20'b00100110110011011010: color_data = 12'b111011101110;
20'b00100110110011011011: color_data = 12'b111011101110;
20'b00100110110011011100: color_data = 12'b111011101110;
20'b00100110110011011101: color_data = 12'b111011101110;
20'b00100110110011011110: color_data = 12'b111011101110;
20'b00100110110011011111: color_data = 12'b111011101110;
20'b00100110110011100000: color_data = 12'b111011101110;
20'b00100110110011100001: color_data = 12'b111011101110;
20'b00100110110011101110: color_data = 12'b111011101110;
20'b00100110110011101111: color_data = 12'b111011101110;
20'b00100110110011110000: color_data = 12'b111011101110;
20'b00100110110011110001: color_data = 12'b111011101110;
20'b00100110110011110010: color_data = 12'b111011101110;
20'b00100110110011110011: color_data = 12'b111011101110;
20'b00100110110011110100: color_data = 12'b111011101110;
20'b00100110110011110101: color_data = 12'b111011101110;
20'b00100110110011110110: color_data = 12'b111011101110;
20'b00100110110011110111: color_data = 12'b111011101110;
20'b00100110110011111001: color_data = 12'b111011101110;
20'b00100110110011111010: color_data = 12'b111011101110;
20'b00100110110011111011: color_data = 12'b111011101110;
20'b00100110110011111100: color_data = 12'b111011101110;
20'b00100110110011111101: color_data = 12'b111011101110;
20'b00100110110011111110: color_data = 12'b111011101110;
20'b00100110110011111111: color_data = 12'b111011101110;
20'b00100110110100000000: color_data = 12'b111011101110;
20'b00100110110100000001: color_data = 12'b111011101110;
20'b00100110110100000010: color_data = 12'b111011101110;
20'b00100110110100100101: color_data = 12'b111011101110;
20'b00100110110100100110: color_data = 12'b111011101110;
20'b00100110110100100111: color_data = 12'b111011101110;
20'b00100110110100101000: color_data = 12'b111011101110;
20'b00100110110100101001: color_data = 12'b111011101110;
20'b00100110110100101010: color_data = 12'b111011101110;
20'b00100110110100101011: color_data = 12'b111011101110;
20'b00100110110100101100: color_data = 12'b111011101110;
20'b00100110110100101101: color_data = 12'b111011101110;
20'b00100110110100101110: color_data = 12'b111011101110;
20'b00100110110100110000: color_data = 12'b111011101110;
20'b00100110110100110001: color_data = 12'b111011101110;
20'b00100110110100110010: color_data = 12'b111011101110;
20'b00100110110100110011: color_data = 12'b111011101110;
20'b00100110110100110100: color_data = 12'b111011101110;
20'b00100110110100110101: color_data = 12'b111011101110;
20'b00100110110100110110: color_data = 12'b111011101110;
20'b00100110110100110111: color_data = 12'b111011101110;
20'b00100110110100111000: color_data = 12'b111011101110;
20'b00100110110100111001: color_data = 12'b111011101110;
20'b00100110110101000110: color_data = 12'b111011101110;
20'b00100110110101000111: color_data = 12'b111011101110;
20'b00100110110101001000: color_data = 12'b111011101110;
20'b00100110110101001001: color_data = 12'b111011101110;
20'b00100110110101001010: color_data = 12'b111011101110;
20'b00100110110101001011: color_data = 12'b111011101110;
20'b00100110110101001100: color_data = 12'b111011101110;
20'b00100110110101001101: color_data = 12'b111011101110;
20'b00100110110101001110: color_data = 12'b111011101110;
20'b00100110110101001111: color_data = 12'b111011101110;
20'b00100110110101010001: color_data = 12'b111011101110;
20'b00100110110101010010: color_data = 12'b111011101110;
20'b00100110110101010011: color_data = 12'b111011101110;
20'b00100110110101010100: color_data = 12'b111011101110;
20'b00100110110101010101: color_data = 12'b111011101110;
20'b00100110110101010110: color_data = 12'b111011101110;
20'b00100110110101010111: color_data = 12'b111011101110;
20'b00100110110101011000: color_data = 12'b111011101110;
20'b00100110110101011001: color_data = 12'b111011101110;
20'b00100110110101011010: color_data = 12'b111011101110;
20'b00100110110101100111: color_data = 12'b111011101110;
20'b00100110110101101000: color_data = 12'b111011101110;
20'b00100110110101101001: color_data = 12'b111011101110;
20'b00100110110101101010: color_data = 12'b111011101110;
20'b00100110110101101011: color_data = 12'b111011101110;
20'b00100110110101101100: color_data = 12'b111011101110;
20'b00100110110101101101: color_data = 12'b111011101110;
20'b00100110110101101110: color_data = 12'b111011101110;
20'b00100110110101101111: color_data = 12'b111011101110;
20'b00100110110101110000: color_data = 12'b111011101110;
20'b00100110110101111101: color_data = 12'b111011101110;
20'b00100110110101111110: color_data = 12'b111011101110;
20'b00100110110101111111: color_data = 12'b111011101110;
20'b00100110110110000000: color_data = 12'b111011101110;
20'b00100110110110000001: color_data = 12'b111011101110;
20'b00100110110110000010: color_data = 12'b111011101110;
20'b00100110110110000011: color_data = 12'b111011101110;
20'b00100110110110000100: color_data = 12'b111011101110;
20'b00100110110110000101: color_data = 12'b111011101110;
20'b00100110110110000110: color_data = 12'b111011101110;
20'b00100110110110001000: color_data = 12'b111011101110;
20'b00100110110110001001: color_data = 12'b111011101110;
20'b00100110110110001010: color_data = 12'b111011101110;
20'b00100110110110001011: color_data = 12'b111011101110;
20'b00100110110110001100: color_data = 12'b111011101110;
20'b00100110110110001101: color_data = 12'b111011101110;
20'b00100110110110001110: color_data = 12'b111011101110;
20'b00100110110110001111: color_data = 12'b111011101110;
20'b00100110110110010000: color_data = 12'b111011101110;
20'b00100110110110010001: color_data = 12'b111011101110;
20'b00100110110110011110: color_data = 12'b111011101110;
20'b00100110110110011111: color_data = 12'b111011101110;
20'b00100110110110100000: color_data = 12'b111011101110;
20'b00100110110110100001: color_data = 12'b111011101110;
20'b00100110110110100010: color_data = 12'b111011101110;
20'b00100110110110100011: color_data = 12'b111011101110;
20'b00100110110110100100: color_data = 12'b111011101110;
20'b00100110110110100101: color_data = 12'b111011101110;
20'b00100110110110100110: color_data = 12'b111011101110;
20'b00100110110110100111: color_data = 12'b111011101110;
20'b00100110110110101001: color_data = 12'b111011101110;
20'b00100110110110101010: color_data = 12'b111011101110;
20'b00100110110110101011: color_data = 12'b111011101110;
20'b00100110110110101100: color_data = 12'b111011101110;
20'b00100110110110101101: color_data = 12'b111011101110;
20'b00100110110110101110: color_data = 12'b111011101110;
20'b00100110110110101111: color_data = 12'b111011101110;
20'b00100110110110110000: color_data = 12'b111011101110;
20'b00100110110110110001: color_data = 12'b111011101110;
20'b00100110110110110010: color_data = 12'b111011101110;
20'b00100110110110110100: color_data = 12'b111011101110;
20'b00100110110110110101: color_data = 12'b111011101110;
20'b00100110110110110110: color_data = 12'b111011101110;
20'b00100110110110110111: color_data = 12'b111011101110;
20'b00100110110110111000: color_data = 12'b111011101110;
20'b00100110110110111001: color_data = 12'b111011101110;
20'b00100110110110111010: color_data = 12'b111011101110;
20'b00100110110110111011: color_data = 12'b111011101110;
20'b00100110110110111100: color_data = 12'b111011101110;
20'b00100110110110111101: color_data = 12'b111011101110;
20'b00100110110110111111: color_data = 12'b111011101110;
20'b00100110110111000000: color_data = 12'b111011101110;
20'b00100110110111000001: color_data = 12'b111011101110;
20'b00100110110111000010: color_data = 12'b111011101110;
20'b00100110110111000011: color_data = 12'b111011101110;
20'b00100110110111000100: color_data = 12'b111011101110;
20'b00100110110111000101: color_data = 12'b111011101110;
20'b00100110110111000110: color_data = 12'b111011101110;
20'b00100110110111000111: color_data = 12'b111011101110;
20'b00100110110111001000: color_data = 12'b111011101110;
20'b00100110110111001010: color_data = 12'b111011101110;
20'b00100110110111001011: color_data = 12'b111011101110;
20'b00100110110111001100: color_data = 12'b111011101110;
20'b00100110110111001101: color_data = 12'b111011101110;
20'b00100110110111001110: color_data = 12'b111011101110;
20'b00100110110111001111: color_data = 12'b111011101110;
20'b00100110110111010000: color_data = 12'b111011101110;
20'b00100110110111010001: color_data = 12'b111011101110;
20'b00100110110111010010: color_data = 12'b111011101110;
20'b00100110110111010011: color_data = 12'b111011101110;
20'b00100111000011000010: color_data = 12'b111011101110;
20'b00100111000011000011: color_data = 12'b111011101110;
20'b00100111000011000100: color_data = 12'b111011101110;
20'b00100111000011000101: color_data = 12'b111011101110;
20'b00100111000011000110: color_data = 12'b111011101110;
20'b00100111000011000111: color_data = 12'b111011101110;
20'b00100111000011001000: color_data = 12'b111011101110;
20'b00100111000011001001: color_data = 12'b111011101110;
20'b00100111000011001010: color_data = 12'b111011101110;
20'b00100111000011001011: color_data = 12'b111011101110;
20'b00100111000011001101: color_data = 12'b111011101110;
20'b00100111000011001110: color_data = 12'b111011101110;
20'b00100111000011001111: color_data = 12'b111011101110;
20'b00100111000011010000: color_data = 12'b111011101110;
20'b00100111000011010001: color_data = 12'b111011101110;
20'b00100111000011010010: color_data = 12'b111011101110;
20'b00100111000011010011: color_data = 12'b111011101110;
20'b00100111000011010100: color_data = 12'b111011101110;
20'b00100111000011010101: color_data = 12'b111011101110;
20'b00100111000011010110: color_data = 12'b111011101110;
20'b00100111000011011000: color_data = 12'b111011101110;
20'b00100111000011011001: color_data = 12'b111011101110;
20'b00100111000011011010: color_data = 12'b111011101110;
20'b00100111000011011011: color_data = 12'b111011101110;
20'b00100111000011011100: color_data = 12'b111011101110;
20'b00100111000011011101: color_data = 12'b111011101110;
20'b00100111000011011110: color_data = 12'b111011101110;
20'b00100111000011011111: color_data = 12'b111011101110;
20'b00100111000011100000: color_data = 12'b111011101110;
20'b00100111000011100001: color_data = 12'b111011101110;
20'b00100111010010010110: color_data = 12'b111011101110;
20'b00100111010010010111: color_data = 12'b111011101110;
20'b00100111010010011000: color_data = 12'b111011101110;
20'b00100111010010011001: color_data = 12'b111011101110;
20'b00100111010010011010: color_data = 12'b111011101110;
20'b00100111010010011011: color_data = 12'b111011101110;
20'b00100111010010011100: color_data = 12'b111011101110;
20'b00100111010010011101: color_data = 12'b111011101110;
20'b00100111010010011110: color_data = 12'b111011101110;
20'b00100111010010011111: color_data = 12'b111011101110;
20'b00100111010010100001: color_data = 12'b111011101110;
20'b00100111010010100010: color_data = 12'b111011101110;
20'b00100111010010100011: color_data = 12'b111011101110;
20'b00100111010010100100: color_data = 12'b111011101110;
20'b00100111010010100101: color_data = 12'b111011101110;
20'b00100111010010100110: color_data = 12'b111011101110;
20'b00100111010010100111: color_data = 12'b111011101110;
20'b00100111010010101000: color_data = 12'b111011101110;
20'b00100111010010101001: color_data = 12'b111011101110;
20'b00100111010010101010: color_data = 12'b111011101110;
20'b00100111010011000010: color_data = 12'b111011101110;
20'b00100111010011000011: color_data = 12'b111011101110;
20'b00100111010011000100: color_data = 12'b111011101110;
20'b00100111010011000101: color_data = 12'b111011101110;
20'b00100111010011000110: color_data = 12'b111011101110;
20'b00100111010011000111: color_data = 12'b111011101110;
20'b00100111010011001000: color_data = 12'b111011101110;
20'b00100111010011001001: color_data = 12'b111011101110;
20'b00100111010011001010: color_data = 12'b111011101110;
20'b00100111010011001011: color_data = 12'b111011101110;
20'b00100111010011001101: color_data = 12'b111011101110;
20'b00100111010011001110: color_data = 12'b111011101110;
20'b00100111010011001111: color_data = 12'b111011101110;
20'b00100111010011010000: color_data = 12'b111011101110;
20'b00100111010011010001: color_data = 12'b111011101110;
20'b00100111010011010010: color_data = 12'b111011101110;
20'b00100111010011010011: color_data = 12'b111011101110;
20'b00100111010011010100: color_data = 12'b111011101110;
20'b00100111010011010101: color_data = 12'b111011101110;
20'b00100111010011010110: color_data = 12'b111011101110;
20'b00100111010011011000: color_data = 12'b111011101110;
20'b00100111010011011001: color_data = 12'b111011101110;
20'b00100111010011011010: color_data = 12'b111011101110;
20'b00100111010011011011: color_data = 12'b111011101110;
20'b00100111010011011100: color_data = 12'b111011101110;
20'b00100111010011011101: color_data = 12'b111011101110;
20'b00100111010011011110: color_data = 12'b111011101110;
20'b00100111010011011111: color_data = 12'b111011101110;
20'b00100111010011100000: color_data = 12'b111011101110;
20'b00100111010011100001: color_data = 12'b111011101110;
20'b00100111010011101110: color_data = 12'b111011101110;
20'b00100111010011101111: color_data = 12'b111011101110;
20'b00100111010011110000: color_data = 12'b111011101110;
20'b00100111010011110001: color_data = 12'b111011101110;
20'b00100111010011110010: color_data = 12'b111011101110;
20'b00100111010011110011: color_data = 12'b111011101110;
20'b00100111010011110100: color_data = 12'b111011101110;
20'b00100111010011110101: color_data = 12'b111011101110;
20'b00100111010011110110: color_data = 12'b111011101110;
20'b00100111010011110111: color_data = 12'b111011101110;
20'b00100111010011111001: color_data = 12'b111011101110;
20'b00100111010011111010: color_data = 12'b111011101110;
20'b00100111010011111011: color_data = 12'b111011101110;
20'b00100111010011111100: color_data = 12'b111011101110;
20'b00100111010011111101: color_data = 12'b111011101110;
20'b00100111010011111110: color_data = 12'b111011101110;
20'b00100111010011111111: color_data = 12'b111011101110;
20'b00100111010100000000: color_data = 12'b111011101110;
20'b00100111010100000001: color_data = 12'b111011101110;
20'b00100111010100000010: color_data = 12'b111011101110;
20'b00100111010100000100: color_data = 12'b111011101110;
20'b00100111010100000101: color_data = 12'b111011101110;
20'b00100111010100000110: color_data = 12'b111011101110;
20'b00100111010100000111: color_data = 12'b111011101110;
20'b00100111010100001000: color_data = 12'b111011101110;
20'b00100111010100001001: color_data = 12'b111011101110;
20'b00100111010100001010: color_data = 12'b111011101110;
20'b00100111010100001011: color_data = 12'b111011101110;
20'b00100111010100001100: color_data = 12'b111011101110;
20'b00100111010100001101: color_data = 12'b111011101110;
20'b00100111010100001111: color_data = 12'b111011101110;
20'b00100111010100010000: color_data = 12'b111011101110;
20'b00100111010100010001: color_data = 12'b111011101110;
20'b00100111010100010010: color_data = 12'b111011101110;
20'b00100111010100010011: color_data = 12'b111011101110;
20'b00100111010100010100: color_data = 12'b111011101110;
20'b00100111010100010101: color_data = 12'b111011101110;
20'b00100111010100010110: color_data = 12'b111011101110;
20'b00100111010100010111: color_data = 12'b111011101110;
20'b00100111010100011000: color_data = 12'b111011101110;
20'b00100111010100011010: color_data = 12'b111011101110;
20'b00100111010100011011: color_data = 12'b111011101110;
20'b00100111010100011100: color_data = 12'b111011101110;
20'b00100111010100011101: color_data = 12'b111011101110;
20'b00100111010100011110: color_data = 12'b111011101110;
20'b00100111010100011111: color_data = 12'b111011101110;
20'b00100111010100100000: color_data = 12'b111011101110;
20'b00100111010100100001: color_data = 12'b111011101110;
20'b00100111010100100010: color_data = 12'b111011101110;
20'b00100111010100100011: color_data = 12'b111011101110;
20'b00100111010100100101: color_data = 12'b111011101110;
20'b00100111010100100110: color_data = 12'b111011101110;
20'b00100111010100100111: color_data = 12'b111011101110;
20'b00100111010100101000: color_data = 12'b111011101110;
20'b00100111010100101001: color_data = 12'b111011101110;
20'b00100111010100101010: color_data = 12'b111011101110;
20'b00100111010100101011: color_data = 12'b111011101110;
20'b00100111010100101100: color_data = 12'b111011101110;
20'b00100111010100101101: color_data = 12'b111011101110;
20'b00100111010100101110: color_data = 12'b111011101110;
20'b00100111010100110000: color_data = 12'b111011101110;
20'b00100111010100110001: color_data = 12'b111011101110;
20'b00100111010100110010: color_data = 12'b111011101110;
20'b00100111010100110011: color_data = 12'b111011101110;
20'b00100111010100110100: color_data = 12'b111011101110;
20'b00100111010100110101: color_data = 12'b111011101110;
20'b00100111010100110110: color_data = 12'b111011101110;
20'b00100111010100110111: color_data = 12'b111011101110;
20'b00100111010100111000: color_data = 12'b111011101110;
20'b00100111010100111001: color_data = 12'b111011101110;
20'b00100111010101000110: color_data = 12'b111011101110;
20'b00100111010101000111: color_data = 12'b111011101110;
20'b00100111010101001000: color_data = 12'b111011101110;
20'b00100111010101001001: color_data = 12'b111011101110;
20'b00100111010101001010: color_data = 12'b111011101110;
20'b00100111010101001011: color_data = 12'b111011101110;
20'b00100111010101001100: color_data = 12'b111011101110;
20'b00100111010101001101: color_data = 12'b111011101110;
20'b00100111010101001110: color_data = 12'b111011101110;
20'b00100111010101001111: color_data = 12'b111011101110;
20'b00100111010101010001: color_data = 12'b111011101110;
20'b00100111010101010010: color_data = 12'b111011101110;
20'b00100111010101010011: color_data = 12'b111011101110;
20'b00100111010101010100: color_data = 12'b111011101110;
20'b00100111010101010101: color_data = 12'b111011101110;
20'b00100111010101010110: color_data = 12'b111011101110;
20'b00100111010101010111: color_data = 12'b111011101110;
20'b00100111010101011000: color_data = 12'b111011101110;
20'b00100111010101011001: color_data = 12'b111011101110;
20'b00100111010101011010: color_data = 12'b111011101110;
20'b00100111010101111101: color_data = 12'b111011101110;
20'b00100111010101111110: color_data = 12'b111011101110;
20'b00100111010101111111: color_data = 12'b111011101110;
20'b00100111010110000000: color_data = 12'b111011101110;
20'b00100111010110000001: color_data = 12'b111011101110;
20'b00100111010110000010: color_data = 12'b111011101110;
20'b00100111010110000011: color_data = 12'b111011101110;
20'b00100111010110000100: color_data = 12'b111011101110;
20'b00100111010110000101: color_data = 12'b111011101110;
20'b00100111010110000110: color_data = 12'b111011101110;
20'b00100111010110001000: color_data = 12'b111011101110;
20'b00100111010110001001: color_data = 12'b111011101110;
20'b00100111010110001010: color_data = 12'b111011101110;
20'b00100111010110001011: color_data = 12'b111011101110;
20'b00100111010110001100: color_data = 12'b111011101110;
20'b00100111010110001101: color_data = 12'b111011101110;
20'b00100111010110001110: color_data = 12'b111011101110;
20'b00100111010110001111: color_data = 12'b111011101110;
20'b00100111010110010000: color_data = 12'b111011101110;
20'b00100111010110010001: color_data = 12'b111011101110;
20'b00100111010110011110: color_data = 12'b111011101110;
20'b00100111010110011111: color_data = 12'b111011101110;
20'b00100111010110100000: color_data = 12'b111011101110;
20'b00100111010110100001: color_data = 12'b111011101110;
20'b00100111010110100010: color_data = 12'b111011101110;
20'b00100111010110100011: color_data = 12'b111011101110;
20'b00100111010110100100: color_data = 12'b111011101110;
20'b00100111010110100101: color_data = 12'b111011101110;
20'b00100111010110100110: color_data = 12'b111011101110;
20'b00100111010110100111: color_data = 12'b111011101110;
20'b00100111010110101001: color_data = 12'b111011101110;
20'b00100111010110101010: color_data = 12'b111011101110;
20'b00100111010110101011: color_data = 12'b111011101110;
20'b00100111010110101100: color_data = 12'b111011101110;
20'b00100111010110101101: color_data = 12'b111011101110;
20'b00100111010110101110: color_data = 12'b111011101110;
20'b00100111010110101111: color_data = 12'b111011101110;
20'b00100111010110110000: color_data = 12'b111011101110;
20'b00100111010110110001: color_data = 12'b111011101110;
20'b00100111010110110010: color_data = 12'b111011101110;
20'b00100111100010010110: color_data = 12'b111011101110;
20'b00100111100010010111: color_data = 12'b111011101110;
20'b00100111100010011000: color_data = 12'b111011101110;
20'b00100111100010011001: color_data = 12'b111011101110;
20'b00100111100010011010: color_data = 12'b111011101110;
20'b00100111100010011011: color_data = 12'b111011101110;
20'b00100111100010011100: color_data = 12'b111011101110;
20'b00100111100010011101: color_data = 12'b111011101110;
20'b00100111100010011110: color_data = 12'b111011101110;
20'b00100111100010011111: color_data = 12'b111011101110;
20'b00100111100010100001: color_data = 12'b111011101110;
20'b00100111100010100010: color_data = 12'b111011101110;
20'b00100111100010100011: color_data = 12'b111011101110;
20'b00100111100010100100: color_data = 12'b111011101110;
20'b00100111100010100101: color_data = 12'b111011101110;
20'b00100111100010100110: color_data = 12'b111011101110;
20'b00100111100010100111: color_data = 12'b111011101110;
20'b00100111100010101000: color_data = 12'b111011101110;
20'b00100111100010101001: color_data = 12'b111011101110;
20'b00100111100010101010: color_data = 12'b111011101110;
20'b00100111100011000010: color_data = 12'b111011101110;
20'b00100111100011000011: color_data = 12'b111011101110;
20'b00100111100011000100: color_data = 12'b111011101110;
20'b00100111100011000101: color_data = 12'b111011101110;
20'b00100111100011000110: color_data = 12'b111011101110;
20'b00100111100011000111: color_data = 12'b111011101110;
20'b00100111100011001000: color_data = 12'b111011101110;
20'b00100111100011001001: color_data = 12'b111011101110;
20'b00100111100011001010: color_data = 12'b111011101110;
20'b00100111100011001011: color_data = 12'b111011101110;
20'b00100111100011001101: color_data = 12'b111011101110;
20'b00100111100011001110: color_data = 12'b111011101110;
20'b00100111100011001111: color_data = 12'b111011101110;
20'b00100111100011010000: color_data = 12'b111011101110;
20'b00100111100011010001: color_data = 12'b111011101110;
20'b00100111100011010010: color_data = 12'b111011101110;
20'b00100111100011010011: color_data = 12'b111011101110;
20'b00100111100011010100: color_data = 12'b111011101110;
20'b00100111100011010101: color_data = 12'b111011101110;
20'b00100111100011010110: color_data = 12'b111011101110;
20'b00100111100011011000: color_data = 12'b111011101110;
20'b00100111100011011001: color_data = 12'b111011101110;
20'b00100111100011011010: color_data = 12'b111011101110;
20'b00100111100011011011: color_data = 12'b111011101110;
20'b00100111100011011100: color_data = 12'b111011101110;
20'b00100111100011011101: color_data = 12'b111011101110;
20'b00100111100011011110: color_data = 12'b111011101110;
20'b00100111100011011111: color_data = 12'b111011101110;
20'b00100111100011100000: color_data = 12'b111011101110;
20'b00100111100011100001: color_data = 12'b111011101110;
20'b00100111100011101110: color_data = 12'b111011101110;
20'b00100111100011101111: color_data = 12'b111011101110;
20'b00100111100011110000: color_data = 12'b111011101110;
20'b00100111100011110001: color_data = 12'b111011101110;
20'b00100111100011110010: color_data = 12'b111011101110;
20'b00100111100011110011: color_data = 12'b111011101110;
20'b00100111100011110100: color_data = 12'b111011101110;
20'b00100111100011110101: color_data = 12'b111011101110;
20'b00100111100011110110: color_data = 12'b111011101110;
20'b00100111100011110111: color_data = 12'b111011101110;
20'b00100111100011111001: color_data = 12'b111011101110;
20'b00100111100011111010: color_data = 12'b111011101110;
20'b00100111100011111011: color_data = 12'b111011101110;
20'b00100111100011111100: color_data = 12'b111011101110;
20'b00100111100011111101: color_data = 12'b111011101110;
20'b00100111100011111110: color_data = 12'b111011101110;
20'b00100111100011111111: color_data = 12'b111011101110;
20'b00100111100100000000: color_data = 12'b111011101110;
20'b00100111100100000001: color_data = 12'b111011101110;
20'b00100111100100000010: color_data = 12'b111011101110;
20'b00100111100100000100: color_data = 12'b111011101110;
20'b00100111100100000101: color_data = 12'b111011101110;
20'b00100111100100000110: color_data = 12'b111011101110;
20'b00100111100100000111: color_data = 12'b111011101110;
20'b00100111100100001000: color_data = 12'b111011101110;
20'b00100111100100001001: color_data = 12'b111011101110;
20'b00100111100100001010: color_data = 12'b111011101110;
20'b00100111100100001011: color_data = 12'b111011101110;
20'b00100111100100001100: color_data = 12'b111011101110;
20'b00100111100100001101: color_data = 12'b111011101110;
20'b00100111100100001111: color_data = 12'b111011101110;
20'b00100111100100010000: color_data = 12'b111011101110;
20'b00100111100100010001: color_data = 12'b111011101110;
20'b00100111100100010010: color_data = 12'b111011101110;
20'b00100111100100010011: color_data = 12'b111011101110;
20'b00100111100100010100: color_data = 12'b111011101110;
20'b00100111100100010101: color_data = 12'b111011101110;
20'b00100111100100010110: color_data = 12'b111011101110;
20'b00100111100100010111: color_data = 12'b111011101110;
20'b00100111100100011000: color_data = 12'b111011101110;
20'b00100111100100011010: color_data = 12'b111011101110;
20'b00100111100100011011: color_data = 12'b111011101110;
20'b00100111100100011100: color_data = 12'b111011101110;
20'b00100111100100011101: color_data = 12'b111011101110;
20'b00100111100100011110: color_data = 12'b111011101110;
20'b00100111100100011111: color_data = 12'b111011101110;
20'b00100111100100100000: color_data = 12'b111011101110;
20'b00100111100100100001: color_data = 12'b111011101110;
20'b00100111100100100010: color_data = 12'b111011101110;
20'b00100111100100100011: color_data = 12'b111011101110;
20'b00100111100100100101: color_data = 12'b111011101110;
20'b00100111100100100110: color_data = 12'b111011101110;
20'b00100111100100100111: color_data = 12'b111011101110;
20'b00100111100100101000: color_data = 12'b111011101110;
20'b00100111100100101001: color_data = 12'b111011101110;
20'b00100111100100101010: color_data = 12'b111011101110;
20'b00100111100100101011: color_data = 12'b111011101110;
20'b00100111100100101100: color_data = 12'b111011101110;
20'b00100111100100101101: color_data = 12'b111011101110;
20'b00100111100100101110: color_data = 12'b111011101110;
20'b00100111100100110000: color_data = 12'b111011101110;
20'b00100111100100110001: color_data = 12'b111011101110;
20'b00100111100100110010: color_data = 12'b111011101110;
20'b00100111100100110011: color_data = 12'b111011101110;
20'b00100111100100110100: color_data = 12'b111011101110;
20'b00100111100100110101: color_data = 12'b111011101110;
20'b00100111100100110110: color_data = 12'b111011101110;
20'b00100111100100110111: color_data = 12'b111011101110;
20'b00100111100100111000: color_data = 12'b111011101110;
20'b00100111100100111001: color_data = 12'b111011101110;
20'b00100111100101000110: color_data = 12'b111011101110;
20'b00100111100101000111: color_data = 12'b111011101110;
20'b00100111100101001000: color_data = 12'b111011101110;
20'b00100111100101001001: color_data = 12'b111011101110;
20'b00100111100101001010: color_data = 12'b111011101110;
20'b00100111100101001011: color_data = 12'b111011101110;
20'b00100111100101001100: color_data = 12'b111011101110;
20'b00100111100101001101: color_data = 12'b111011101110;
20'b00100111100101001110: color_data = 12'b111011101110;
20'b00100111100101001111: color_data = 12'b111011101110;
20'b00100111100101010001: color_data = 12'b111011101110;
20'b00100111100101010010: color_data = 12'b111011101110;
20'b00100111100101010011: color_data = 12'b111011101110;
20'b00100111100101010100: color_data = 12'b111011101110;
20'b00100111100101010101: color_data = 12'b111011101110;
20'b00100111100101010110: color_data = 12'b111011101110;
20'b00100111100101010111: color_data = 12'b111011101110;
20'b00100111100101011000: color_data = 12'b111011101110;
20'b00100111100101011001: color_data = 12'b111011101110;
20'b00100111100101011010: color_data = 12'b111011101110;
20'b00100111100101111101: color_data = 12'b111011101110;
20'b00100111100101111110: color_data = 12'b111011101110;
20'b00100111100101111111: color_data = 12'b111011101110;
20'b00100111100110000000: color_data = 12'b111011101110;
20'b00100111100110000001: color_data = 12'b111011101110;
20'b00100111100110000010: color_data = 12'b111011101110;
20'b00100111100110000011: color_data = 12'b111011101110;
20'b00100111100110000100: color_data = 12'b111011101110;
20'b00100111100110000101: color_data = 12'b111011101110;
20'b00100111100110000110: color_data = 12'b111011101110;
20'b00100111100110001000: color_data = 12'b111011101110;
20'b00100111100110001001: color_data = 12'b111011101110;
20'b00100111100110001010: color_data = 12'b111011101110;
20'b00100111100110001011: color_data = 12'b111011101110;
20'b00100111100110001100: color_data = 12'b111011101110;
20'b00100111100110001101: color_data = 12'b111011101110;
20'b00100111100110001110: color_data = 12'b111011101110;
20'b00100111100110001111: color_data = 12'b111011101110;
20'b00100111100110010000: color_data = 12'b111011101110;
20'b00100111100110010001: color_data = 12'b111011101110;
20'b00100111100110011110: color_data = 12'b111011101110;
20'b00100111100110011111: color_data = 12'b111011101110;
20'b00100111100110100000: color_data = 12'b111011101110;
20'b00100111100110100001: color_data = 12'b111011101110;
20'b00100111100110100010: color_data = 12'b111011101110;
20'b00100111100110100011: color_data = 12'b111011101110;
20'b00100111100110100100: color_data = 12'b111011101110;
20'b00100111100110100101: color_data = 12'b111011101110;
20'b00100111100110100110: color_data = 12'b111011101110;
20'b00100111100110100111: color_data = 12'b111011101110;
20'b00100111100110101001: color_data = 12'b111011101110;
20'b00100111100110101010: color_data = 12'b111011101110;
20'b00100111100110101011: color_data = 12'b111011101110;
20'b00100111100110101100: color_data = 12'b111011101110;
20'b00100111100110101101: color_data = 12'b111011101110;
20'b00100111100110101110: color_data = 12'b111011101110;
20'b00100111100110101111: color_data = 12'b111011101110;
20'b00100111100110110000: color_data = 12'b111011101110;
20'b00100111100110110001: color_data = 12'b111011101110;
20'b00100111100110110010: color_data = 12'b111011101110;
20'b00100111110010010110: color_data = 12'b111011101110;
20'b00100111110010010111: color_data = 12'b111011101110;
20'b00100111110010011000: color_data = 12'b111011101110;
20'b00100111110010011001: color_data = 12'b111011101110;
20'b00100111110010011010: color_data = 12'b111011101110;
20'b00100111110010011011: color_data = 12'b111011101110;
20'b00100111110010011100: color_data = 12'b111011101110;
20'b00100111110010011101: color_data = 12'b111011101110;
20'b00100111110010011110: color_data = 12'b111011101110;
20'b00100111110010011111: color_data = 12'b111011101110;
20'b00100111110010100001: color_data = 12'b111011101110;
20'b00100111110010100010: color_data = 12'b111011101110;
20'b00100111110010100011: color_data = 12'b111011101110;
20'b00100111110010100100: color_data = 12'b111011101110;
20'b00100111110010100101: color_data = 12'b111011101110;
20'b00100111110010100110: color_data = 12'b111011101110;
20'b00100111110010100111: color_data = 12'b111011101110;
20'b00100111110010101000: color_data = 12'b111011101110;
20'b00100111110010101001: color_data = 12'b111011101110;
20'b00100111110010101010: color_data = 12'b111011101110;
20'b00100111110011000010: color_data = 12'b111011101110;
20'b00100111110011000011: color_data = 12'b111011101110;
20'b00100111110011000100: color_data = 12'b111011101110;
20'b00100111110011000101: color_data = 12'b111011101110;
20'b00100111110011000110: color_data = 12'b111011101110;
20'b00100111110011000111: color_data = 12'b111011101110;
20'b00100111110011001000: color_data = 12'b111011101110;
20'b00100111110011001001: color_data = 12'b111011101110;
20'b00100111110011001010: color_data = 12'b111011101110;
20'b00100111110011001011: color_data = 12'b111011101110;
20'b00100111110011001101: color_data = 12'b111011101110;
20'b00100111110011001110: color_data = 12'b111011101110;
20'b00100111110011001111: color_data = 12'b111011101110;
20'b00100111110011010000: color_data = 12'b111011101110;
20'b00100111110011010001: color_data = 12'b111011101110;
20'b00100111110011010010: color_data = 12'b111011101110;
20'b00100111110011010011: color_data = 12'b111011101110;
20'b00100111110011010100: color_data = 12'b111011101110;
20'b00100111110011010101: color_data = 12'b111011101110;
20'b00100111110011010110: color_data = 12'b111011101110;
20'b00100111110011011000: color_data = 12'b111011101110;
20'b00100111110011011001: color_data = 12'b111011101110;
20'b00100111110011011010: color_data = 12'b111011101110;
20'b00100111110011011011: color_data = 12'b111011101110;
20'b00100111110011011100: color_data = 12'b111011101110;
20'b00100111110011011101: color_data = 12'b111011101110;
20'b00100111110011011110: color_data = 12'b111011101110;
20'b00100111110011011111: color_data = 12'b111011101110;
20'b00100111110011100000: color_data = 12'b111011101110;
20'b00100111110011100001: color_data = 12'b111011101110;
20'b00100111110011101110: color_data = 12'b111011101110;
20'b00100111110011101111: color_data = 12'b111011101110;
20'b00100111110011110000: color_data = 12'b111011101110;
20'b00100111110011110001: color_data = 12'b111011101110;
20'b00100111110011110010: color_data = 12'b111011101110;
20'b00100111110011110011: color_data = 12'b111011101110;
20'b00100111110011110100: color_data = 12'b111011101110;
20'b00100111110011110101: color_data = 12'b111011101110;
20'b00100111110011110110: color_data = 12'b111011101110;
20'b00100111110011110111: color_data = 12'b111011101110;
20'b00100111110011111001: color_data = 12'b111011101110;
20'b00100111110011111010: color_data = 12'b111011101110;
20'b00100111110011111011: color_data = 12'b111011101110;
20'b00100111110011111100: color_data = 12'b111011101110;
20'b00100111110011111101: color_data = 12'b111011101110;
20'b00100111110011111110: color_data = 12'b111011101110;
20'b00100111110011111111: color_data = 12'b111011101110;
20'b00100111110100000000: color_data = 12'b111011101110;
20'b00100111110100000001: color_data = 12'b111011101110;
20'b00100111110100000010: color_data = 12'b111011101110;
20'b00100111110100000100: color_data = 12'b111011101110;
20'b00100111110100000101: color_data = 12'b111011101110;
20'b00100111110100000110: color_data = 12'b111011101110;
20'b00100111110100000111: color_data = 12'b111011101110;
20'b00100111110100001000: color_data = 12'b111011101110;
20'b00100111110100001001: color_data = 12'b111011101110;
20'b00100111110100001010: color_data = 12'b111011101110;
20'b00100111110100001011: color_data = 12'b111011101110;
20'b00100111110100001100: color_data = 12'b111011101110;
20'b00100111110100001101: color_data = 12'b111011101110;
20'b00100111110100001111: color_data = 12'b111011101110;
20'b00100111110100010000: color_data = 12'b111011101110;
20'b00100111110100010001: color_data = 12'b111011101110;
20'b00100111110100010010: color_data = 12'b111011101110;
20'b00100111110100010011: color_data = 12'b111011101110;
20'b00100111110100010100: color_data = 12'b111011101110;
20'b00100111110100010101: color_data = 12'b111011101110;
20'b00100111110100010110: color_data = 12'b111011101110;
20'b00100111110100010111: color_data = 12'b111011101110;
20'b00100111110100011000: color_data = 12'b111011101110;
20'b00100111110100011010: color_data = 12'b111011101110;
20'b00100111110100011011: color_data = 12'b111011101110;
20'b00100111110100011100: color_data = 12'b111011101110;
20'b00100111110100011101: color_data = 12'b111011101110;
20'b00100111110100011110: color_data = 12'b111011101110;
20'b00100111110100011111: color_data = 12'b111011101110;
20'b00100111110100100000: color_data = 12'b111011101110;
20'b00100111110100100001: color_data = 12'b111011101110;
20'b00100111110100100010: color_data = 12'b111011101110;
20'b00100111110100100011: color_data = 12'b111011101110;
20'b00100111110100100101: color_data = 12'b111011101110;
20'b00100111110100100110: color_data = 12'b111011101110;
20'b00100111110100100111: color_data = 12'b111011101110;
20'b00100111110100101000: color_data = 12'b111011101110;
20'b00100111110100101001: color_data = 12'b111011101110;
20'b00100111110100101010: color_data = 12'b111011101110;
20'b00100111110100101011: color_data = 12'b111011101110;
20'b00100111110100101100: color_data = 12'b111011101110;
20'b00100111110100101101: color_data = 12'b111011101110;
20'b00100111110100101110: color_data = 12'b111011101110;
20'b00100111110100110000: color_data = 12'b111011101110;
20'b00100111110100110001: color_data = 12'b111011101110;
20'b00100111110100110010: color_data = 12'b111011101110;
20'b00100111110100110011: color_data = 12'b111011101110;
20'b00100111110100110100: color_data = 12'b111011101110;
20'b00100111110100110101: color_data = 12'b111011101110;
20'b00100111110100110110: color_data = 12'b111011101110;
20'b00100111110100110111: color_data = 12'b111011101110;
20'b00100111110100111000: color_data = 12'b111011101110;
20'b00100111110100111001: color_data = 12'b111011101110;
20'b00100111110101000110: color_data = 12'b111011101110;
20'b00100111110101000111: color_data = 12'b111011101110;
20'b00100111110101001000: color_data = 12'b111011101110;
20'b00100111110101001001: color_data = 12'b111011101110;
20'b00100111110101001010: color_data = 12'b111011101110;
20'b00100111110101001011: color_data = 12'b111011101110;
20'b00100111110101001100: color_data = 12'b111011101110;
20'b00100111110101001101: color_data = 12'b111011101110;
20'b00100111110101001110: color_data = 12'b111011101110;
20'b00100111110101001111: color_data = 12'b111011101110;
20'b00100111110101010001: color_data = 12'b111011101110;
20'b00100111110101010010: color_data = 12'b111011101110;
20'b00100111110101010011: color_data = 12'b111011101110;
20'b00100111110101010100: color_data = 12'b111011101110;
20'b00100111110101010101: color_data = 12'b111011101110;
20'b00100111110101010110: color_data = 12'b111011101110;
20'b00100111110101010111: color_data = 12'b111011101110;
20'b00100111110101011000: color_data = 12'b111011101110;
20'b00100111110101011001: color_data = 12'b111011101110;
20'b00100111110101011010: color_data = 12'b111011101110;
20'b00100111110101111101: color_data = 12'b111011101110;
20'b00100111110101111110: color_data = 12'b111011101110;
20'b00100111110101111111: color_data = 12'b111011101110;
20'b00100111110110000000: color_data = 12'b111011101110;
20'b00100111110110000001: color_data = 12'b111011101110;
20'b00100111110110000010: color_data = 12'b111011101110;
20'b00100111110110000011: color_data = 12'b111011101110;
20'b00100111110110000100: color_data = 12'b111011101110;
20'b00100111110110000101: color_data = 12'b111011101110;
20'b00100111110110000110: color_data = 12'b111011101110;
20'b00100111110110001000: color_data = 12'b111011101110;
20'b00100111110110001001: color_data = 12'b111011101110;
20'b00100111110110001010: color_data = 12'b111011101110;
20'b00100111110110001011: color_data = 12'b111011101110;
20'b00100111110110001100: color_data = 12'b111011101110;
20'b00100111110110001101: color_data = 12'b111011101110;
20'b00100111110110001110: color_data = 12'b111011101110;
20'b00100111110110001111: color_data = 12'b111011101110;
20'b00100111110110010000: color_data = 12'b111011101110;
20'b00100111110110010001: color_data = 12'b111011101110;
20'b00100111110110011110: color_data = 12'b111011101110;
20'b00100111110110011111: color_data = 12'b111011101110;
20'b00100111110110100000: color_data = 12'b111011101110;
20'b00100111110110100001: color_data = 12'b111011101110;
20'b00100111110110100010: color_data = 12'b111011101110;
20'b00100111110110100011: color_data = 12'b111011101110;
20'b00100111110110100100: color_data = 12'b111011101110;
20'b00100111110110100101: color_data = 12'b111011101110;
20'b00100111110110100110: color_data = 12'b111011101110;
20'b00100111110110100111: color_data = 12'b111011101110;
20'b00100111110110101001: color_data = 12'b111011101110;
20'b00100111110110101010: color_data = 12'b111011101110;
20'b00100111110110101011: color_data = 12'b111011101110;
20'b00100111110110101100: color_data = 12'b111011101110;
20'b00100111110110101101: color_data = 12'b111011101110;
20'b00100111110110101110: color_data = 12'b111011101110;
20'b00100111110110101111: color_data = 12'b111011101110;
20'b00100111110110110000: color_data = 12'b111011101110;
20'b00100111110110110001: color_data = 12'b111011101110;
20'b00100111110110110010: color_data = 12'b111011101110;
20'b00101000000010010110: color_data = 12'b111011101110;
20'b00101000000010010111: color_data = 12'b111011101110;
20'b00101000000010011000: color_data = 12'b111011101110;
20'b00101000000010011001: color_data = 12'b111011101110;
20'b00101000000010011010: color_data = 12'b111011101110;
20'b00101000000010011011: color_data = 12'b111011101110;
20'b00101000000010011100: color_data = 12'b111011101110;
20'b00101000000010011101: color_data = 12'b111011101110;
20'b00101000000010011110: color_data = 12'b111011101110;
20'b00101000000010011111: color_data = 12'b111011101110;
20'b00101000000010100001: color_data = 12'b111011101110;
20'b00101000000010100010: color_data = 12'b111011101110;
20'b00101000000010100011: color_data = 12'b111011101110;
20'b00101000000010100100: color_data = 12'b111011101110;
20'b00101000000010100101: color_data = 12'b111011101110;
20'b00101000000010100110: color_data = 12'b111011101110;
20'b00101000000010100111: color_data = 12'b111011101110;
20'b00101000000010101000: color_data = 12'b111011101110;
20'b00101000000010101001: color_data = 12'b111011101110;
20'b00101000000010101010: color_data = 12'b111011101110;
20'b00101000000011000010: color_data = 12'b111011101110;
20'b00101000000011000011: color_data = 12'b111011101110;
20'b00101000000011000100: color_data = 12'b111011101110;
20'b00101000000011000101: color_data = 12'b111011101110;
20'b00101000000011000110: color_data = 12'b111011101110;
20'b00101000000011000111: color_data = 12'b111011101110;
20'b00101000000011001000: color_data = 12'b111011101110;
20'b00101000000011001001: color_data = 12'b111011101110;
20'b00101000000011001010: color_data = 12'b111011101110;
20'b00101000000011001011: color_data = 12'b111011101110;
20'b00101000000011001101: color_data = 12'b111011101110;
20'b00101000000011001110: color_data = 12'b111011101110;
20'b00101000000011001111: color_data = 12'b111011101110;
20'b00101000000011010000: color_data = 12'b111011101110;
20'b00101000000011010001: color_data = 12'b111011101110;
20'b00101000000011010010: color_data = 12'b111011101110;
20'b00101000000011010011: color_data = 12'b111011101110;
20'b00101000000011010100: color_data = 12'b111011101110;
20'b00101000000011010101: color_data = 12'b111011101110;
20'b00101000000011010110: color_data = 12'b111011101110;
20'b00101000000011011000: color_data = 12'b111011101110;
20'b00101000000011011001: color_data = 12'b111011101110;
20'b00101000000011011010: color_data = 12'b111011101110;
20'b00101000000011011011: color_data = 12'b111011101110;
20'b00101000000011011100: color_data = 12'b111011101110;
20'b00101000000011011101: color_data = 12'b111011101110;
20'b00101000000011011110: color_data = 12'b111011101110;
20'b00101000000011011111: color_data = 12'b111011101110;
20'b00101000000011100000: color_data = 12'b111011101110;
20'b00101000000011100001: color_data = 12'b111011101110;
20'b00101000000011101110: color_data = 12'b111011101110;
20'b00101000000011101111: color_data = 12'b111011101110;
20'b00101000000011110000: color_data = 12'b111011101110;
20'b00101000000011110001: color_data = 12'b111011101110;
20'b00101000000011110010: color_data = 12'b111011101110;
20'b00101000000011110011: color_data = 12'b111011101110;
20'b00101000000011110100: color_data = 12'b111011101110;
20'b00101000000011110101: color_data = 12'b111011101110;
20'b00101000000011110110: color_data = 12'b111011101110;
20'b00101000000011110111: color_data = 12'b111011101110;
20'b00101000000011111001: color_data = 12'b111011101110;
20'b00101000000011111010: color_data = 12'b111011101110;
20'b00101000000011111011: color_data = 12'b111011101110;
20'b00101000000011111100: color_data = 12'b111011101110;
20'b00101000000011111101: color_data = 12'b111011101110;
20'b00101000000011111110: color_data = 12'b111011101110;
20'b00101000000011111111: color_data = 12'b111011101110;
20'b00101000000100000000: color_data = 12'b111011101110;
20'b00101000000100000001: color_data = 12'b111011101110;
20'b00101000000100000010: color_data = 12'b111011101110;
20'b00101000000100000100: color_data = 12'b111011101110;
20'b00101000000100000101: color_data = 12'b111011101110;
20'b00101000000100000110: color_data = 12'b111011101110;
20'b00101000000100000111: color_data = 12'b111011101110;
20'b00101000000100001000: color_data = 12'b111011101110;
20'b00101000000100001001: color_data = 12'b111011101110;
20'b00101000000100001010: color_data = 12'b111011101110;
20'b00101000000100001011: color_data = 12'b111011101110;
20'b00101000000100001100: color_data = 12'b111011101110;
20'b00101000000100001101: color_data = 12'b111011101110;
20'b00101000000100001111: color_data = 12'b111011101110;
20'b00101000000100010000: color_data = 12'b111011101110;
20'b00101000000100010001: color_data = 12'b111011101110;
20'b00101000000100010010: color_data = 12'b111011101110;
20'b00101000000100010011: color_data = 12'b111011101110;
20'b00101000000100010100: color_data = 12'b111011101110;
20'b00101000000100010101: color_data = 12'b111011101110;
20'b00101000000100010110: color_data = 12'b111011101110;
20'b00101000000100010111: color_data = 12'b111011101110;
20'b00101000000100011000: color_data = 12'b111011101110;
20'b00101000000100011010: color_data = 12'b111011101110;
20'b00101000000100011011: color_data = 12'b111011101110;
20'b00101000000100011100: color_data = 12'b111011101110;
20'b00101000000100011101: color_data = 12'b111011101110;
20'b00101000000100011110: color_data = 12'b111011101110;
20'b00101000000100011111: color_data = 12'b111011101110;
20'b00101000000100100000: color_data = 12'b111011101110;
20'b00101000000100100001: color_data = 12'b111011101110;
20'b00101000000100100010: color_data = 12'b111011101110;
20'b00101000000100100011: color_data = 12'b111011101110;
20'b00101000000100100101: color_data = 12'b111011101110;
20'b00101000000100100110: color_data = 12'b111011101110;
20'b00101000000100100111: color_data = 12'b111011101110;
20'b00101000000100101000: color_data = 12'b111011101110;
20'b00101000000100101001: color_data = 12'b111011101110;
20'b00101000000100101010: color_data = 12'b111011101110;
20'b00101000000100101011: color_data = 12'b111011101110;
20'b00101000000100101100: color_data = 12'b111011101110;
20'b00101000000100101101: color_data = 12'b111011101110;
20'b00101000000100101110: color_data = 12'b111011101110;
20'b00101000000100110000: color_data = 12'b111011101110;
20'b00101000000100110001: color_data = 12'b111011101110;
20'b00101000000100110010: color_data = 12'b111011101110;
20'b00101000000100110011: color_data = 12'b111011101110;
20'b00101000000100110100: color_data = 12'b111011101110;
20'b00101000000100110101: color_data = 12'b111011101110;
20'b00101000000100110110: color_data = 12'b111011101110;
20'b00101000000100110111: color_data = 12'b111011101110;
20'b00101000000100111000: color_data = 12'b111011101110;
20'b00101000000100111001: color_data = 12'b111011101110;
20'b00101000000101000110: color_data = 12'b111011101110;
20'b00101000000101000111: color_data = 12'b111011101110;
20'b00101000000101001000: color_data = 12'b111011101110;
20'b00101000000101001001: color_data = 12'b111011101110;
20'b00101000000101001010: color_data = 12'b111011101110;
20'b00101000000101001011: color_data = 12'b111011101110;
20'b00101000000101001100: color_data = 12'b111011101110;
20'b00101000000101001101: color_data = 12'b111011101110;
20'b00101000000101001110: color_data = 12'b111011101110;
20'b00101000000101001111: color_data = 12'b111011101110;
20'b00101000000101010001: color_data = 12'b111011101110;
20'b00101000000101010010: color_data = 12'b111011101110;
20'b00101000000101010011: color_data = 12'b111011101110;
20'b00101000000101010100: color_data = 12'b111011101110;
20'b00101000000101010101: color_data = 12'b111011101110;
20'b00101000000101010110: color_data = 12'b111011101110;
20'b00101000000101010111: color_data = 12'b111011101110;
20'b00101000000101011000: color_data = 12'b111011101110;
20'b00101000000101011001: color_data = 12'b111011101110;
20'b00101000000101011010: color_data = 12'b111011101110;
20'b00101000000101111101: color_data = 12'b111011101110;
20'b00101000000101111110: color_data = 12'b111011101110;
20'b00101000000101111111: color_data = 12'b111011101110;
20'b00101000000110000000: color_data = 12'b111011101110;
20'b00101000000110000001: color_data = 12'b111011101110;
20'b00101000000110000010: color_data = 12'b111011101110;
20'b00101000000110000011: color_data = 12'b111011101110;
20'b00101000000110000100: color_data = 12'b111011101110;
20'b00101000000110000101: color_data = 12'b111011101110;
20'b00101000000110000110: color_data = 12'b111011101110;
20'b00101000000110001000: color_data = 12'b111011101110;
20'b00101000000110001001: color_data = 12'b111011101110;
20'b00101000000110001010: color_data = 12'b111011101110;
20'b00101000000110001011: color_data = 12'b111011101110;
20'b00101000000110001100: color_data = 12'b111011101110;
20'b00101000000110001101: color_data = 12'b111011101110;
20'b00101000000110001110: color_data = 12'b111011101110;
20'b00101000000110001111: color_data = 12'b111011101110;
20'b00101000000110010000: color_data = 12'b111011101110;
20'b00101000000110010001: color_data = 12'b111011101110;
20'b00101000000110011110: color_data = 12'b111011101110;
20'b00101000000110011111: color_data = 12'b111011101110;
20'b00101000000110100000: color_data = 12'b111011101110;
20'b00101000000110100001: color_data = 12'b111011101110;
20'b00101000000110100010: color_data = 12'b111011101110;
20'b00101000000110100011: color_data = 12'b111011101110;
20'b00101000000110100100: color_data = 12'b111011101110;
20'b00101000000110100101: color_data = 12'b111011101110;
20'b00101000000110100110: color_data = 12'b111011101110;
20'b00101000000110100111: color_data = 12'b111011101110;
20'b00101000000110101001: color_data = 12'b111011101110;
20'b00101000000110101010: color_data = 12'b111011101110;
20'b00101000000110101011: color_data = 12'b111011101110;
20'b00101000000110101100: color_data = 12'b111011101110;
20'b00101000000110101101: color_data = 12'b111011101110;
20'b00101000000110101110: color_data = 12'b111011101110;
20'b00101000000110101111: color_data = 12'b111011101110;
20'b00101000000110110000: color_data = 12'b111011101110;
20'b00101000000110110001: color_data = 12'b111011101110;
20'b00101000000110110010: color_data = 12'b111011101110;
20'b00101000010010010110: color_data = 12'b111011101110;
20'b00101000010010010111: color_data = 12'b111011101110;
20'b00101000010010011000: color_data = 12'b111011101110;
20'b00101000010010011001: color_data = 12'b111011101110;
20'b00101000010010011010: color_data = 12'b111011101110;
20'b00101000010010011011: color_data = 12'b111011101110;
20'b00101000010010011100: color_data = 12'b111011101110;
20'b00101000010010011101: color_data = 12'b111011101110;
20'b00101000010010011110: color_data = 12'b111011101110;
20'b00101000010010011111: color_data = 12'b111011101110;
20'b00101000010010100001: color_data = 12'b111011101110;
20'b00101000010010100010: color_data = 12'b111011101110;
20'b00101000010010100011: color_data = 12'b111011101110;
20'b00101000010010100100: color_data = 12'b111011101110;
20'b00101000010010100101: color_data = 12'b111011101110;
20'b00101000010010100110: color_data = 12'b111011101110;
20'b00101000010010100111: color_data = 12'b111011101110;
20'b00101000010010101000: color_data = 12'b111011101110;
20'b00101000010010101001: color_data = 12'b111011101110;
20'b00101000010010101010: color_data = 12'b111011101110;
20'b00101000010011000010: color_data = 12'b111011101110;
20'b00101000010011000011: color_data = 12'b111011101110;
20'b00101000010011000100: color_data = 12'b111011101110;
20'b00101000010011000101: color_data = 12'b111011101110;
20'b00101000010011000110: color_data = 12'b111011101110;
20'b00101000010011000111: color_data = 12'b111011101110;
20'b00101000010011001000: color_data = 12'b111011101110;
20'b00101000010011001001: color_data = 12'b111011101110;
20'b00101000010011001010: color_data = 12'b111011101110;
20'b00101000010011001011: color_data = 12'b111011101110;
20'b00101000010011001101: color_data = 12'b111011101110;
20'b00101000010011001110: color_data = 12'b111011101110;
20'b00101000010011001111: color_data = 12'b111011101110;
20'b00101000010011010000: color_data = 12'b111011101110;
20'b00101000010011010001: color_data = 12'b111011101110;
20'b00101000010011010010: color_data = 12'b111011101110;
20'b00101000010011010011: color_data = 12'b111011101110;
20'b00101000010011010100: color_data = 12'b111011101110;
20'b00101000010011010101: color_data = 12'b111011101110;
20'b00101000010011010110: color_data = 12'b111011101110;
20'b00101000010011011000: color_data = 12'b111011101110;
20'b00101000010011011001: color_data = 12'b111011101110;
20'b00101000010011011010: color_data = 12'b111011101110;
20'b00101000010011011011: color_data = 12'b111011101110;
20'b00101000010011011100: color_data = 12'b111011101110;
20'b00101000010011011101: color_data = 12'b111011101110;
20'b00101000010011011110: color_data = 12'b111011101110;
20'b00101000010011011111: color_data = 12'b111011101110;
20'b00101000010011100000: color_data = 12'b111011101110;
20'b00101000010011100001: color_data = 12'b111011101110;
20'b00101000010011101110: color_data = 12'b111011101110;
20'b00101000010011101111: color_data = 12'b111011101110;
20'b00101000010011110000: color_data = 12'b111011101110;
20'b00101000010011110001: color_data = 12'b111011101110;
20'b00101000010011110010: color_data = 12'b111011101110;
20'b00101000010011110011: color_data = 12'b111011101110;
20'b00101000010011110100: color_data = 12'b111011101110;
20'b00101000010011110101: color_data = 12'b111011101110;
20'b00101000010011110110: color_data = 12'b111011101110;
20'b00101000010011110111: color_data = 12'b111011101110;
20'b00101000010011111001: color_data = 12'b111011101110;
20'b00101000010011111010: color_data = 12'b111011101110;
20'b00101000010011111011: color_data = 12'b111011101110;
20'b00101000010011111100: color_data = 12'b111011101110;
20'b00101000010011111101: color_data = 12'b111011101110;
20'b00101000010011111110: color_data = 12'b111011101110;
20'b00101000010011111111: color_data = 12'b111011101110;
20'b00101000010100000000: color_data = 12'b111011101110;
20'b00101000010100000001: color_data = 12'b111011101110;
20'b00101000010100000010: color_data = 12'b111011101110;
20'b00101000010100000100: color_data = 12'b111011101110;
20'b00101000010100000101: color_data = 12'b111011101110;
20'b00101000010100000110: color_data = 12'b111011101110;
20'b00101000010100000111: color_data = 12'b111011101110;
20'b00101000010100001000: color_data = 12'b111011101110;
20'b00101000010100001001: color_data = 12'b111011101110;
20'b00101000010100001010: color_data = 12'b111011101110;
20'b00101000010100001011: color_data = 12'b111011101110;
20'b00101000010100001100: color_data = 12'b111011101110;
20'b00101000010100001101: color_data = 12'b111011101110;
20'b00101000010100001111: color_data = 12'b111011101110;
20'b00101000010100010000: color_data = 12'b111011101110;
20'b00101000010100010001: color_data = 12'b111011101110;
20'b00101000010100010010: color_data = 12'b111011101110;
20'b00101000010100010011: color_data = 12'b111011101110;
20'b00101000010100010100: color_data = 12'b111011101110;
20'b00101000010100010101: color_data = 12'b111011101110;
20'b00101000010100010110: color_data = 12'b111011101110;
20'b00101000010100010111: color_data = 12'b111011101110;
20'b00101000010100011000: color_data = 12'b111011101110;
20'b00101000010100011010: color_data = 12'b111011101110;
20'b00101000010100011011: color_data = 12'b111011101110;
20'b00101000010100011100: color_data = 12'b111011101110;
20'b00101000010100011101: color_data = 12'b111011101110;
20'b00101000010100011110: color_data = 12'b111011101110;
20'b00101000010100011111: color_data = 12'b111011101110;
20'b00101000010100100000: color_data = 12'b111011101110;
20'b00101000010100100001: color_data = 12'b111011101110;
20'b00101000010100100010: color_data = 12'b111011101110;
20'b00101000010100100011: color_data = 12'b111011101110;
20'b00101000010100100101: color_data = 12'b111011101110;
20'b00101000010100100110: color_data = 12'b111011101110;
20'b00101000010100100111: color_data = 12'b111011101110;
20'b00101000010100101000: color_data = 12'b111011101110;
20'b00101000010100101001: color_data = 12'b111011101110;
20'b00101000010100101010: color_data = 12'b111011101110;
20'b00101000010100101011: color_data = 12'b111011101110;
20'b00101000010100101100: color_data = 12'b111011101110;
20'b00101000010100101101: color_data = 12'b111011101110;
20'b00101000010100101110: color_data = 12'b111011101110;
20'b00101000010100110000: color_data = 12'b111011101110;
20'b00101000010100110001: color_data = 12'b111011101110;
20'b00101000010100110010: color_data = 12'b111011101110;
20'b00101000010100110011: color_data = 12'b111011101110;
20'b00101000010100110100: color_data = 12'b111011101110;
20'b00101000010100110101: color_data = 12'b111011101110;
20'b00101000010100110110: color_data = 12'b111011101110;
20'b00101000010100110111: color_data = 12'b111011101110;
20'b00101000010100111000: color_data = 12'b111011101110;
20'b00101000010100111001: color_data = 12'b111011101110;
20'b00101000010101000110: color_data = 12'b111011101110;
20'b00101000010101000111: color_data = 12'b111011101110;
20'b00101000010101001000: color_data = 12'b111011101110;
20'b00101000010101001001: color_data = 12'b111011101110;
20'b00101000010101001010: color_data = 12'b111011101110;
20'b00101000010101001011: color_data = 12'b111011101110;
20'b00101000010101001100: color_data = 12'b111011101110;
20'b00101000010101001101: color_data = 12'b111011101110;
20'b00101000010101001110: color_data = 12'b111011101110;
20'b00101000010101001111: color_data = 12'b111011101110;
20'b00101000010101010001: color_data = 12'b111011101110;
20'b00101000010101010010: color_data = 12'b111011101110;
20'b00101000010101010011: color_data = 12'b111011101110;
20'b00101000010101010100: color_data = 12'b111011101110;
20'b00101000010101010101: color_data = 12'b111011101110;
20'b00101000010101010110: color_data = 12'b111011101110;
20'b00101000010101010111: color_data = 12'b111011101110;
20'b00101000010101011000: color_data = 12'b111011101110;
20'b00101000010101011001: color_data = 12'b111011101110;
20'b00101000010101011010: color_data = 12'b111011101110;
20'b00101000010101111101: color_data = 12'b111011101110;
20'b00101000010101111110: color_data = 12'b111011101110;
20'b00101000010101111111: color_data = 12'b111011101110;
20'b00101000010110000000: color_data = 12'b111011101110;
20'b00101000010110000001: color_data = 12'b111011101110;
20'b00101000010110000010: color_data = 12'b111011101110;
20'b00101000010110000011: color_data = 12'b111011101110;
20'b00101000010110000100: color_data = 12'b111011101110;
20'b00101000010110000101: color_data = 12'b111011101110;
20'b00101000010110000110: color_data = 12'b111011101110;
20'b00101000010110001000: color_data = 12'b111011101110;
20'b00101000010110001001: color_data = 12'b111011101110;
20'b00101000010110001010: color_data = 12'b111011101110;
20'b00101000010110001011: color_data = 12'b111011101110;
20'b00101000010110001100: color_data = 12'b111011101110;
20'b00101000010110001101: color_data = 12'b111011101110;
20'b00101000010110001110: color_data = 12'b111011101110;
20'b00101000010110001111: color_data = 12'b111011101110;
20'b00101000010110010000: color_data = 12'b111011101110;
20'b00101000010110010001: color_data = 12'b111011101110;
20'b00101000010110011110: color_data = 12'b111011101110;
20'b00101000010110011111: color_data = 12'b111011101110;
20'b00101000010110100000: color_data = 12'b111011101110;
20'b00101000010110100001: color_data = 12'b111011101110;
20'b00101000010110100010: color_data = 12'b111011101110;
20'b00101000010110100011: color_data = 12'b111011101110;
20'b00101000010110100100: color_data = 12'b111011101110;
20'b00101000010110100101: color_data = 12'b111011101110;
20'b00101000010110100110: color_data = 12'b111011101110;
20'b00101000010110100111: color_data = 12'b111011101110;
20'b00101000010110101001: color_data = 12'b111011101110;
20'b00101000010110101010: color_data = 12'b111011101110;
20'b00101000010110101011: color_data = 12'b111011101110;
20'b00101000010110101100: color_data = 12'b111011101110;
20'b00101000010110101101: color_data = 12'b111011101110;
20'b00101000010110101110: color_data = 12'b111011101110;
20'b00101000010110101111: color_data = 12'b111011101110;
20'b00101000010110110000: color_data = 12'b111011101110;
20'b00101000010110110001: color_data = 12'b111011101110;
20'b00101000010110110010: color_data = 12'b111011101110;
20'b00101000100010010110: color_data = 12'b111011101110;
20'b00101000100010010111: color_data = 12'b111011101110;
20'b00101000100010011000: color_data = 12'b111011101110;
20'b00101000100010011001: color_data = 12'b111011101110;
20'b00101000100010011010: color_data = 12'b111011101110;
20'b00101000100010011011: color_data = 12'b111011101110;
20'b00101000100010011100: color_data = 12'b111011101110;
20'b00101000100010011101: color_data = 12'b111011101110;
20'b00101000100010011110: color_data = 12'b111011101110;
20'b00101000100010011111: color_data = 12'b111011101110;
20'b00101000100010100001: color_data = 12'b111011101110;
20'b00101000100010100010: color_data = 12'b111011101110;
20'b00101000100010100011: color_data = 12'b111011101110;
20'b00101000100010100100: color_data = 12'b111011101110;
20'b00101000100010100101: color_data = 12'b111011101110;
20'b00101000100010100110: color_data = 12'b111011101110;
20'b00101000100010100111: color_data = 12'b111011101110;
20'b00101000100010101000: color_data = 12'b111011101110;
20'b00101000100010101001: color_data = 12'b111011101110;
20'b00101000100010101010: color_data = 12'b111011101110;
20'b00101000100011000010: color_data = 12'b111011101110;
20'b00101000100011000011: color_data = 12'b111011101110;
20'b00101000100011000100: color_data = 12'b111011101110;
20'b00101000100011000101: color_data = 12'b111011101110;
20'b00101000100011000110: color_data = 12'b111011101110;
20'b00101000100011000111: color_data = 12'b111011101110;
20'b00101000100011001000: color_data = 12'b111011101110;
20'b00101000100011001001: color_data = 12'b111011101110;
20'b00101000100011001010: color_data = 12'b111011101110;
20'b00101000100011001011: color_data = 12'b111011101110;
20'b00101000100011001101: color_data = 12'b111011101110;
20'b00101000100011001110: color_data = 12'b111011101110;
20'b00101000100011001111: color_data = 12'b111011101110;
20'b00101000100011010000: color_data = 12'b111011101110;
20'b00101000100011010001: color_data = 12'b111011101110;
20'b00101000100011010010: color_data = 12'b111011101110;
20'b00101000100011010011: color_data = 12'b111011101110;
20'b00101000100011010100: color_data = 12'b111011101110;
20'b00101000100011010101: color_data = 12'b111011101110;
20'b00101000100011010110: color_data = 12'b111011101110;
20'b00101000100011011000: color_data = 12'b111011101110;
20'b00101000100011011001: color_data = 12'b111011101110;
20'b00101000100011011010: color_data = 12'b111011101110;
20'b00101000100011011011: color_data = 12'b111011101110;
20'b00101000100011011100: color_data = 12'b111011101110;
20'b00101000100011011101: color_data = 12'b111011101110;
20'b00101000100011011110: color_data = 12'b111011101110;
20'b00101000100011011111: color_data = 12'b111011101110;
20'b00101000100011100000: color_data = 12'b111011101110;
20'b00101000100011100001: color_data = 12'b111011101110;
20'b00101000100011101110: color_data = 12'b111011101110;
20'b00101000100011101111: color_data = 12'b111011101110;
20'b00101000100011110000: color_data = 12'b111011101110;
20'b00101000100011110001: color_data = 12'b111011101110;
20'b00101000100011110010: color_data = 12'b111011101110;
20'b00101000100011110011: color_data = 12'b111011101110;
20'b00101000100011110100: color_data = 12'b111011101110;
20'b00101000100011110101: color_data = 12'b111011101110;
20'b00101000100011110110: color_data = 12'b111011101110;
20'b00101000100011110111: color_data = 12'b111011101110;
20'b00101000100011111001: color_data = 12'b111011101110;
20'b00101000100011111010: color_data = 12'b111011101110;
20'b00101000100011111011: color_data = 12'b111011101110;
20'b00101000100011111100: color_data = 12'b111011101110;
20'b00101000100011111101: color_data = 12'b111011101110;
20'b00101000100011111110: color_data = 12'b111011101110;
20'b00101000100011111111: color_data = 12'b111011101110;
20'b00101000100100000000: color_data = 12'b111011101110;
20'b00101000100100000001: color_data = 12'b111011101110;
20'b00101000100100000010: color_data = 12'b111011101110;
20'b00101000100100000100: color_data = 12'b111011101110;
20'b00101000100100000101: color_data = 12'b111011101110;
20'b00101000100100000110: color_data = 12'b111011101110;
20'b00101000100100000111: color_data = 12'b111011101110;
20'b00101000100100001000: color_data = 12'b111011101110;
20'b00101000100100001001: color_data = 12'b111011101110;
20'b00101000100100001010: color_data = 12'b111011101110;
20'b00101000100100001011: color_data = 12'b111011101110;
20'b00101000100100001100: color_data = 12'b111011101110;
20'b00101000100100001101: color_data = 12'b111011101110;
20'b00101000100100001111: color_data = 12'b111011101110;
20'b00101000100100010000: color_data = 12'b111011101110;
20'b00101000100100010001: color_data = 12'b111011101110;
20'b00101000100100010010: color_data = 12'b111011101110;
20'b00101000100100010011: color_data = 12'b111011101110;
20'b00101000100100010100: color_data = 12'b111011101110;
20'b00101000100100010101: color_data = 12'b111011101110;
20'b00101000100100010110: color_data = 12'b111011101110;
20'b00101000100100010111: color_data = 12'b111011101110;
20'b00101000100100011000: color_data = 12'b111011101110;
20'b00101000100100011010: color_data = 12'b111011101110;
20'b00101000100100011011: color_data = 12'b111011101110;
20'b00101000100100011100: color_data = 12'b111011101110;
20'b00101000100100011101: color_data = 12'b111011101110;
20'b00101000100100011110: color_data = 12'b111011101110;
20'b00101000100100011111: color_data = 12'b111011101110;
20'b00101000100100100000: color_data = 12'b111011101110;
20'b00101000100100100001: color_data = 12'b111011101110;
20'b00101000100100100010: color_data = 12'b111011101110;
20'b00101000100100100011: color_data = 12'b111011101110;
20'b00101000100100100101: color_data = 12'b111011101110;
20'b00101000100100100110: color_data = 12'b111011101110;
20'b00101000100100100111: color_data = 12'b111011101110;
20'b00101000100100101000: color_data = 12'b111011101110;
20'b00101000100100101001: color_data = 12'b111011101110;
20'b00101000100100101010: color_data = 12'b111011101110;
20'b00101000100100101011: color_data = 12'b111011101110;
20'b00101000100100101100: color_data = 12'b111011101110;
20'b00101000100100101101: color_data = 12'b111011101110;
20'b00101000100100101110: color_data = 12'b111011101110;
20'b00101000100100110000: color_data = 12'b111011101110;
20'b00101000100100110001: color_data = 12'b111011101110;
20'b00101000100100110010: color_data = 12'b111011101110;
20'b00101000100100110011: color_data = 12'b111011101110;
20'b00101000100100110100: color_data = 12'b111011101110;
20'b00101000100100110101: color_data = 12'b111011101110;
20'b00101000100100110110: color_data = 12'b111011101110;
20'b00101000100100110111: color_data = 12'b111011101110;
20'b00101000100100111000: color_data = 12'b111011101110;
20'b00101000100100111001: color_data = 12'b111011101110;
20'b00101000100101000110: color_data = 12'b111011101110;
20'b00101000100101000111: color_data = 12'b111011101110;
20'b00101000100101001000: color_data = 12'b111011101110;
20'b00101000100101001001: color_data = 12'b111011101110;
20'b00101000100101001010: color_data = 12'b111011101110;
20'b00101000100101001011: color_data = 12'b111011101110;
20'b00101000100101001100: color_data = 12'b111011101110;
20'b00101000100101001101: color_data = 12'b111011101110;
20'b00101000100101001110: color_data = 12'b111011101110;
20'b00101000100101001111: color_data = 12'b111011101110;
20'b00101000100101010001: color_data = 12'b111011101110;
20'b00101000100101010010: color_data = 12'b111011101110;
20'b00101000100101010011: color_data = 12'b111011101110;
20'b00101000100101010100: color_data = 12'b111011101110;
20'b00101000100101010101: color_data = 12'b111011101110;
20'b00101000100101010110: color_data = 12'b111011101110;
20'b00101000100101010111: color_data = 12'b111011101110;
20'b00101000100101011000: color_data = 12'b111011101110;
20'b00101000100101011001: color_data = 12'b111011101110;
20'b00101000100101011010: color_data = 12'b111011101110;
20'b00101000100101111101: color_data = 12'b111011101110;
20'b00101000100101111110: color_data = 12'b111011101110;
20'b00101000100101111111: color_data = 12'b111011101110;
20'b00101000100110000000: color_data = 12'b111011101110;
20'b00101000100110000001: color_data = 12'b111011101110;
20'b00101000100110000010: color_data = 12'b111011101110;
20'b00101000100110000011: color_data = 12'b111011101110;
20'b00101000100110000100: color_data = 12'b111011101110;
20'b00101000100110000101: color_data = 12'b111011101110;
20'b00101000100110000110: color_data = 12'b111011101110;
20'b00101000100110001000: color_data = 12'b111011101110;
20'b00101000100110001001: color_data = 12'b111011101110;
20'b00101000100110001010: color_data = 12'b111011101110;
20'b00101000100110001011: color_data = 12'b111011101110;
20'b00101000100110001100: color_data = 12'b111011101110;
20'b00101000100110001101: color_data = 12'b111011101110;
20'b00101000100110001110: color_data = 12'b111011101110;
20'b00101000100110001111: color_data = 12'b111011101110;
20'b00101000100110010000: color_data = 12'b111011101110;
20'b00101000100110010001: color_data = 12'b111011101110;
20'b00101000100110011110: color_data = 12'b111011101110;
20'b00101000100110011111: color_data = 12'b111011101110;
20'b00101000100110100000: color_data = 12'b111011101110;
20'b00101000100110100001: color_data = 12'b111011101110;
20'b00101000100110100010: color_data = 12'b111011101110;
20'b00101000100110100011: color_data = 12'b111011101110;
20'b00101000100110100100: color_data = 12'b111011101110;
20'b00101000100110100101: color_data = 12'b111011101110;
20'b00101000100110100110: color_data = 12'b111011101110;
20'b00101000100110100111: color_data = 12'b111011101110;
20'b00101000100110101001: color_data = 12'b111011101110;
20'b00101000100110101010: color_data = 12'b111011101110;
20'b00101000100110101011: color_data = 12'b111011101110;
20'b00101000100110101100: color_data = 12'b111011101110;
20'b00101000100110101101: color_data = 12'b111011101110;
20'b00101000100110101110: color_data = 12'b111011101110;
20'b00101000100110101111: color_data = 12'b111011101110;
20'b00101000100110110000: color_data = 12'b111011101110;
20'b00101000100110110001: color_data = 12'b111011101110;
20'b00101000100110110010: color_data = 12'b111011101110;
20'b00101000110010010110: color_data = 12'b111011101110;
20'b00101000110010010111: color_data = 12'b111011101110;
20'b00101000110010011000: color_data = 12'b111011101110;
20'b00101000110010011001: color_data = 12'b111011101110;
20'b00101000110010011010: color_data = 12'b111011101110;
20'b00101000110010011011: color_data = 12'b111011101110;
20'b00101000110010011100: color_data = 12'b111011101110;
20'b00101000110010011101: color_data = 12'b111011101110;
20'b00101000110010011110: color_data = 12'b111011101110;
20'b00101000110010011111: color_data = 12'b111011101110;
20'b00101000110010100001: color_data = 12'b111011101110;
20'b00101000110010100010: color_data = 12'b111011101110;
20'b00101000110010100011: color_data = 12'b111011101110;
20'b00101000110010100100: color_data = 12'b111011101110;
20'b00101000110010100101: color_data = 12'b111011101110;
20'b00101000110010100110: color_data = 12'b111011101110;
20'b00101000110010100111: color_data = 12'b111011101110;
20'b00101000110010101000: color_data = 12'b111011101110;
20'b00101000110010101001: color_data = 12'b111011101110;
20'b00101000110010101010: color_data = 12'b111011101110;
20'b00101000110011000010: color_data = 12'b111011101110;
20'b00101000110011000011: color_data = 12'b111011101110;
20'b00101000110011000100: color_data = 12'b111011101110;
20'b00101000110011000101: color_data = 12'b111011101110;
20'b00101000110011000110: color_data = 12'b111011101110;
20'b00101000110011000111: color_data = 12'b111011101110;
20'b00101000110011001000: color_data = 12'b111011101110;
20'b00101000110011001001: color_data = 12'b111011101110;
20'b00101000110011001010: color_data = 12'b111011101110;
20'b00101000110011001011: color_data = 12'b111011101110;
20'b00101000110011001101: color_data = 12'b111011101110;
20'b00101000110011001110: color_data = 12'b111011101110;
20'b00101000110011001111: color_data = 12'b111011101110;
20'b00101000110011010000: color_data = 12'b111011101110;
20'b00101000110011010001: color_data = 12'b111011101110;
20'b00101000110011010010: color_data = 12'b111011101110;
20'b00101000110011010011: color_data = 12'b111011101110;
20'b00101000110011010100: color_data = 12'b111011101110;
20'b00101000110011010101: color_data = 12'b111011101110;
20'b00101000110011010110: color_data = 12'b111011101110;
20'b00101000110011011000: color_data = 12'b111011101110;
20'b00101000110011011001: color_data = 12'b111011101110;
20'b00101000110011011010: color_data = 12'b111011101110;
20'b00101000110011011011: color_data = 12'b111011101110;
20'b00101000110011011100: color_data = 12'b111011101110;
20'b00101000110011011101: color_data = 12'b111011101110;
20'b00101000110011011110: color_data = 12'b111011101110;
20'b00101000110011011111: color_data = 12'b111011101110;
20'b00101000110011100000: color_data = 12'b111011101110;
20'b00101000110011100001: color_data = 12'b111011101110;
20'b00101000110011101110: color_data = 12'b111011101110;
20'b00101000110011101111: color_data = 12'b111011101110;
20'b00101000110011110000: color_data = 12'b111011101110;
20'b00101000110011110001: color_data = 12'b111011101110;
20'b00101000110011110010: color_data = 12'b111011101110;
20'b00101000110011110011: color_data = 12'b111011101110;
20'b00101000110011110100: color_data = 12'b111011101110;
20'b00101000110011110101: color_data = 12'b111011101110;
20'b00101000110011110110: color_data = 12'b111011101110;
20'b00101000110011110111: color_data = 12'b111011101110;
20'b00101000110011111001: color_data = 12'b111011101110;
20'b00101000110011111010: color_data = 12'b111011101110;
20'b00101000110011111011: color_data = 12'b111011101110;
20'b00101000110011111100: color_data = 12'b111011101110;
20'b00101000110011111101: color_data = 12'b111011101110;
20'b00101000110011111110: color_data = 12'b111011101110;
20'b00101000110011111111: color_data = 12'b111011101110;
20'b00101000110100000000: color_data = 12'b111011101110;
20'b00101000110100000001: color_data = 12'b111011101110;
20'b00101000110100000010: color_data = 12'b111011101110;
20'b00101000110100000100: color_data = 12'b111011101110;
20'b00101000110100000101: color_data = 12'b111011101110;
20'b00101000110100000110: color_data = 12'b111011101110;
20'b00101000110100000111: color_data = 12'b111011101110;
20'b00101000110100001000: color_data = 12'b111011101110;
20'b00101000110100001001: color_data = 12'b111011101110;
20'b00101000110100001010: color_data = 12'b111011101110;
20'b00101000110100001011: color_data = 12'b111011101110;
20'b00101000110100001100: color_data = 12'b111011101110;
20'b00101000110100001101: color_data = 12'b111011101110;
20'b00101000110100001111: color_data = 12'b111011101110;
20'b00101000110100010000: color_data = 12'b111011101110;
20'b00101000110100010001: color_data = 12'b111011101110;
20'b00101000110100010010: color_data = 12'b111011101110;
20'b00101000110100010011: color_data = 12'b111011101110;
20'b00101000110100010100: color_data = 12'b111011101110;
20'b00101000110100010101: color_data = 12'b111011101110;
20'b00101000110100010110: color_data = 12'b111011101110;
20'b00101000110100010111: color_data = 12'b111011101110;
20'b00101000110100011000: color_data = 12'b111011101110;
20'b00101000110100011010: color_data = 12'b111011101110;
20'b00101000110100011011: color_data = 12'b111011101110;
20'b00101000110100011100: color_data = 12'b111011101110;
20'b00101000110100011101: color_data = 12'b111011101110;
20'b00101000110100011110: color_data = 12'b111011101110;
20'b00101000110100011111: color_data = 12'b111011101110;
20'b00101000110100100000: color_data = 12'b111011101110;
20'b00101000110100100001: color_data = 12'b111011101110;
20'b00101000110100100010: color_data = 12'b111011101110;
20'b00101000110100100011: color_data = 12'b111011101110;
20'b00101000110100100101: color_data = 12'b111011101110;
20'b00101000110100100110: color_data = 12'b111011101110;
20'b00101000110100100111: color_data = 12'b111011101110;
20'b00101000110100101000: color_data = 12'b111011101110;
20'b00101000110100101001: color_data = 12'b111011101110;
20'b00101000110100101010: color_data = 12'b111011101110;
20'b00101000110100101011: color_data = 12'b111011101110;
20'b00101000110100101100: color_data = 12'b111011101110;
20'b00101000110100101101: color_data = 12'b111011101110;
20'b00101000110100101110: color_data = 12'b111011101110;
20'b00101000110100110000: color_data = 12'b111011101110;
20'b00101000110100110001: color_data = 12'b111011101110;
20'b00101000110100110010: color_data = 12'b111011101110;
20'b00101000110100110011: color_data = 12'b111011101110;
20'b00101000110100110100: color_data = 12'b111011101110;
20'b00101000110100110101: color_data = 12'b111011101110;
20'b00101000110100110110: color_data = 12'b111011101110;
20'b00101000110100110111: color_data = 12'b111011101110;
20'b00101000110100111000: color_data = 12'b111011101110;
20'b00101000110100111001: color_data = 12'b111011101110;
20'b00101000110101000110: color_data = 12'b111011101110;
20'b00101000110101000111: color_data = 12'b111011101110;
20'b00101000110101001000: color_data = 12'b111011101110;
20'b00101000110101001001: color_data = 12'b111011101110;
20'b00101000110101001010: color_data = 12'b111011101110;
20'b00101000110101001011: color_data = 12'b111011101110;
20'b00101000110101001100: color_data = 12'b111011101110;
20'b00101000110101001101: color_data = 12'b111011101110;
20'b00101000110101001110: color_data = 12'b111011101110;
20'b00101000110101001111: color_data = 12'b111011101110;
20'b00101000110101010001: color_data = 12'b111011101110;
20'b00101000110101010010: color_data = 12'b111011101110;
20'b00101000110101010011: color_data = 12'b111011101110;
20'b00101000110101010100: color_data = 12'b111011101110;
20'b00101000110101010101: color_data = 12'b111011101110;
20'b00101000110101010110: color_data = 12'b111011101110;
20'b00101000110101010111: color_data = 12'b111011101110;
20'b00101000110101011000: color_data = 12'b111011101110;
20'b00101000110101011001: color_data = 12'b111011101110;
20'b00101000110101011010: color_data = 12'b111011101110;
20'b00101000110101111101: color_data = 12'b111011101110;
20'b00101000110101111110: color_data = 12'b111011101110;
20'b00101000110101111111: color_data = 12'b111011101110;
20'b00101000110110000000: color_data = 12'b111011101110;
20'b00101000110110000001: color_data = 12'b111011101110;
20'b00101000110110000010: color_data = 12'b111011101110;
20'b00101000110110000011: color_data = 12'b111011101110;
20'b00101000110110000100: color_data = 12'b111011101110;
20'b00101000110110000101: color_data = 12'b111011101110;
20'b00101000110110000110: color_data = 12'b111011101110;
20'b00101000110110001000: color_data = 12'b111011101110;
20'b00101000110110001001: color_data = 12'b111011101110;
20'b00101000110110001010: color_data = 12'b111011101110;
20'b00101000110110001011: color_data = 12'b111011101110;
20'b00101000110110001100: color_data = 12'b111011101110;
20'b00101000110110001101: color_data = 12'b111011101110;
20'b00101000110110001110: color_data = 12'b111011101110;
20'b00101000110110001111: color_data = 12'b111011101110;
20'b00101000110110010000: color_data = 12'b111011101110;
20'b00101000110110010001: color_data = 12'b111011101110;
20'b00101000110110011110: color_data = 12'b111011101110;
20'b00101000110110011111: color_data = 12'b111011101110;
20'b00101000110110100000: color_data = 12'b111011101110;
20'b00101000110110100001: color_data = 12'b111011101110;
20'b00101000110110100010: color_data = 12'b111011101110;
20'b00101000110110100011: color_data = 12'b111011101110;
20'b00101000110110100100: color_data = 12'b111011101110;
20'b00101000110110100101: color_data = 12'b111011101110;
20'b00101000110110100110: color_data = 12'b111011101110;
20'b00101000110110100111: color_data = 12'b111011101110;
20'b00101000110110101001: color_data = 12'b111011101110;
20'b00101000110110101010: color_data = 12'b111011101110;
20'b00101000110110101011: color_data = 12'b111011101110;
20'b00101000110110101100: color_data = 12'b111011101110;
20'b00101000110110101101: color_data = 12'b111011101110;
20'b00101000110110101110: color_data = 12'b111011101110;
20'b00101000110110101111: color_data = 12'b111011101110;
20'b00101000110110110000: color_data = 12'b111011101110;
20'b00101000110110110001: color_data = 12'b111011101110;
20'b00101000110110110010: color_data = 12'b111011101110;
20'b00101001000010010110: color_data = 12'b111011101110;
20'b00101001000010010111: color_data = 12'b111011101110;
20'b00101001000010011000: color_data = 12'b111011101110;
20'b00101001000010011001: color_data = 12'b111011101110;
20'b00101001000010011010: color_data = 12'b111011101110;
20'b00101001000010011011: color_data = 12'b111011101110;
20'b00101001000010011100: color_data = 12'b111011101110;
20'b00101001000010011101: color_data = 12'b111011101110;
20'b00101001000010011110: color_data = 12'b111011101110;
20'b00101001000010011111: color_data = 12'b111011101110;
20'b00101001000010100001: color_data = 12'b111011101110;
20'b00101001000010100010: color_data = 12'b111011101110;
20'b00101001000010100011: color_data = 12'b111011101110;
20'b00101001000010100100: color_data = 12'b111011101110;
20'b00101001000010100101: color_data = 12'b111011101110;
20'b00101001000010100110: color_data = 12'b111011101110;
20'b00101001000010100111: color_data = 12'b111011101110;
20'b00101001000010101000: color_data = 12'b111011101110;
20'b00101001000010101001: color_data = 12'b111011101110;
20'b00101001000010101010: color_data = 12'b111011101110;
20'b00101001000011000010: color_data = 12'b111011101110;
20'b00101001000011000011: color_data = 12'b111011101110;
20'b00101001000011000100: color_data = 12'b111011101110;
20'b00101001000011000101: color_data = 12'b111011101110;
20'b00101001000011000110: color_data = 12'b111011101110;
20'b00101001000011000111: color_data = 12'b111011101110;
20'b00101001000011001000: color_data = 12'b111011101110;
20'b00101001000011001001: color_data = 12'b111011101110;
20'b00101001000011001010: color_data = 12'b111011101110;
20'b00101001000011001011: color_data = 12'b111011101110;
20'b00101001000011001101: color_data = 12'b111011101110;
20'b00101001000011001110: color_data = 12'b111011101110;
20'b00101001000011001111: color_data = 12'b111011101110;
20'b00101001000011010000: color_data = 12'b111011101110;
20'b00101001000011010001: color_data = 12'b111011101110;
20'b00101001000011010010: color_data = 12'b111011101110;
20'b00101001000011010011: color_data = 12'b111011101110;
20'b00101001000011010100: color_data = 12'b111011101110;
20'b00101001000011010101: color_data = 12'b111011101110;
20'b00101001000011010110: color_data = 12'b111011101110;
20'b00101001000011011000: color_data = 12'b111011101110;
20'b00101001000011011001: color_data = 12'b111011101110;
20'b00101001000011011010: color_data = 12'b111011101110;
20'b00101001000011011011: color_data = 12'b111011101110;
20'b00101001000011011100: color_data = 12'b111011101110;
20'b00101001000011011101: color_data = 12'b111011101110;
20'b00101001000011011110: color_data = 12'b111011101110;
20'b00101001000011011111: color_data = 12'b111011101110;
20'b00101001000011100000: color_data = 12'b111011101110;
20'b00101001000011100001: color_data = 12'b111011101110;
20'b00101001000011101110: color_data = 12'b111011101110;
20'b00101001000011101111: color_data = 12'b111011101110;
20'b00101001000011110000: color_data = 12'b111011101110;
20'b00101001000011110001: color_data = 12'b111011101110;
20'b00101001000011110010: color_data = 12'b111011101110;
20'b00101001000011110011: color_data = 12'b111011101110;
20'b00101001000011110100: color_data = 12'b111011101110;
20'b00101001000011110101: color_data = 12'b111011101110;
20'b00101001000011110110: color_data = 12'b111011101110;
20'b00101001000011110111: color_data = 12'b111011101110;
20'b00101001000011111001: color_data = 12'b111011101110;
20'b00101001000011111010: color_data = 12'b111011101110;
20'b00101001000011111011: color_data = 12'b111011101110;
20'b00101001000011111100: color_data = 12'b111011101110;
20'b00101001000011111101: color_data = 12'b111011101110;
20'b00101001000011111110: color_data = 12'b111011101110;
20'b00101001000011111111: color_data = 12'b111011101110;
20'b00101001000100000000: color_data = 12'b111011101110;
20'b00101001000100000001: color_data = 12'b111011101110;
20'b00101001000100000010: color_data = 12'b111011101110;
20'b00101001000100000100: color_data = 12'b111011101110;
20'b00101001000100000101: color_data = 12'b111011101110;
20'b00101001000100000110: color_data = 12'b111011101110;
20'b00101001000100000111: color_data = 12'b111011101110;
20'b00101001000100001000: color_data = 12'b111011101110;
20'b00101001000100001001: color_data = 12'b111011101110;
20'b00101001000100001010: color_data = 12'b111011101110;
20'b00101001000100001011: color_data = 12'b111011101110;
20'b00101001000100001100: color_data = 12'b111011101110;
20'b00101001000100001101: color_data = 12'b111011101110;
20'b00101001000100001111: color_data = 12'b111011101110;
20'b00101001000100010000: color_data = 12'b111011101110;
20'b00101001000100010001: color_data = 12'b111011101110;
20'b00101001000100010010: color_data = 12'b111011101110;
20'b00101001000100010011: color_data = 12'b111011101110;
20'b00101001000100010100: color_data = 12'b111011101110;
20'b00101001000100010101: color_data = 12'b111011101110;
20'b00101001000100010110: color_data = 12'b111011101110;
20'b00101001000100010111: color_data = 12'b111011101110;
20'b00101001000100011000: color_data = 12'b111011101110;
20'b00101001000100011010: color_data = 12'b111011101110;
20'b00101001000100011011: color_data = 12'b111011101110;
20'b00101001000100011100: color_data = 12'b111011101110;
20'b00101001000100011101: color_data = 12'b111011101110;
20'b00101001000100011110: color_data = 12'b111011101110;
20'b00101001000100011111: color_data = 12'b111011101110;
20'b00101001000100100000: color_data = 12'b111011101110;
20'b00101001000100100001: color_data = 12'b111011101110;
20'b00101001000100100010: color_data = 12'b111011101110;
20'b00101001000100100011: color_data = 12'b111011101110;
20'b00101001000100100101: color_data = 12'b111011101110;
20'b00101001000100100110: color_data = 12'b111011101110;
20'b00101001000100100111: color_data = 12'b111011101110;
20'b00101001000100101000: color_data = 12'b111011101110;
20'b00101001000100101001: color_data = 12'b111011101110;
20'b00101001000100101010: color_data = 12'b111011101110;
20'b00101001000100101011: color_data = 12'b111011101110;
20'b00101001000100101100: color_data = 12'b111011101110;
20'b00101001000100101101: color_data = 12'b111011101110;
20'b00101001000100101110: color_data = 12'b111011101110;
20'b00101001000100110000: color_data = 12'b111011101110;
20'b00101001000100110001: color_data = 12'b111011101110;
20'b00101001000100110010: color_data = 12'b111011101110;
20'b00101001000100110011: color_data = 12'b111011101110;
20'b00101001000100110100: color_data = 12'b111011101110;
20'b00101001000100110101: color_data = 12'b111011101110;
20'b00101001000100110110: color_data = 12'b111011101110;
20'b00101001000100110111: color_data = 12'b111011101110;
20'b00101001000100111000: color_data = 12'b111011101110;
20'b00101001000100111001: color_data = 12'b111011101110;
20'b00101001000101000110: color_data = 12'b111011101110;
20'b00101001000101000111: color_data = 12'b111011101110;
20'b00101001000101001000: color_data = 12'b111011101110;
20'b00101001000101001001: color_data = 12'b111011101110;
20'b00101001000101001010: color_data = 12'b111011101110;
20'b00101001000101001011: color_data = 12'b111011101110;
20'b00101001000101001100: color_data = 12'b111011101110;
20'b00101001000101001101: color_data = 12'b111011101110;
20'b00101001000101001110: color_data = 12'b111011101110;
20'b00101001000101001111: color_data = 12'b111011101110;
20'b00101001000101010001: color_data = 12'b111011101110;
20'b00101001000101010010: color_data = 12'b111011101110;
20'b00101001000101010011: color_data = 12'b111011101110;
20'b00101001000101010100: color_data = 12'b111011101110;
20'b00101001000101010101: color_data = 12'b111011101110;
20'b00101001000101010110: color_data = 12'b111011101110;
20'b00101001000101010111: color_data = 12'b111011101110;
20'b00101001000101011000: color_data = 12'b111011101110;
20'b00101001000101011001: color_data = 12'b111011101110;
20'b00101001000101011010: color_data = 12'b111011101110;
20'b00101001000101111101: color_data = 12'b111011101110;
20'b00101001000101111110: color_data = 12'b111011101110;
20'b00101001000101111111: color_data = 12'b111011101110;
20'b00101001000110000000: color_data = 12'b111011101110;
20'b00101001000110000001: color_data = 12'b111011101110;
20'b00101001000110000010: color_data = 12'b111011101110;
20'b00101001000110000011: color_data = 12'b111011101110;
20'b00101001000110000100: color_data = 12'b111011101110;
20'b00101001000110000101: color_data = 12'b111011101110;
20'b00101001000110000110: color_data = 12'b111011101110;
20'b00101001000110001000: color_data = 12'b111011101110;
20'b00101001000110001001: color_data = 12'b111011101110;
20'b00101001000110001010: color_data = 12'b111011101110;
20'b00101001000110001011: color_data = 12'b111011101110;
20'b00101001000110001100: color_data = 12'b111011101110;
20'b00101001000110001101: color_data = 12'b111011101110;
20'b00101001000110001110: color_data = 12'b111011101110;
20'b00101001000110001111: color_data = 12'b111011101110;
20'b00101001000110010000: color_data = 12'b111011101110;
20'b00101001000110010001: color_data = 12'b111011101110;
20'b00101001000110011110: color_data = 12'b111011101110;
20'b00101001000110011111: color_data = 12'b111011101110;
20'b00101001000110100000: color_data = 12'b111011101110;
20'b00101001000110100001: color_data = 12'b111011101110;
20'b00101001000110100010: color_data = 12'b111011101110;
20'b00101001000110100011: color_data = 12'b111011101110;
20'b00101001000110100100: color_data = 12'b111011101110;
20'b00101001000110100101: color_data = 12'b111011101110;
20'b00101001000110100110: color_data = 12'b111011101110;
20'b00101001000110100111: color_data = 12'b111011101110;
20'b00101001000110101001: color_data = 12'b111011101110;
20'b00101001000110101010: color_data = 12'b111011101110;
20'b00101001000110101011: color_data = 12'b111011101110;
20'b00101001000110101100: color_data = 12'b111011101110;
20'b00101001000110101101: color_data = 12'b111011101110;
20'b00101001000110101110: color_data = 12'b111011101110;
20'b00101001000110101111: color_data = 12'b111011101110;
20'b00101001000110110000: color_data = 12'b111011101110;
20'b00101001000110110001: color_data = 12'b111011101110;
20'b00101001000110110010: color_data = 12'b111011101110;
20'b00101001010010010110: color_data = 12'b111011101110;
20'b00101001010010010111: color_data = 12'b111011101110;
20'b00101001010010011000: color_data = 12'b111011101110;
20'b00101001010010011001: color_data = 12'b111011101110;
20'b00101001010010011010: color_data = 12'b111011101110;
20'b00101001010010011011: color_data = 12'b111011101110;
20'b00101001010010011100: color_data = 12'b111011101110;
20'b00101001010010011101: color_data = 12'b111011101110;
20'b00101001010010011110: color_data = 12'b111011101110;
20'b00101001010010011111: color_data = 12'b111011101110;
20'b00101001010010100001: color_data = 12'b111011101110;
20'b00101001010010100010: color_data = 12'b111011101110;
20'b00101001010010100011: color_data = 12'b111011101110;
20'b00101001010010100100: color_data = 12'b111011101110;
20'b00101001010010100101: color_data = 12'b111011101110;
20'b00101001010010100110: color_data = 12'b111011101110;
20'b00101001010010100111: color_data = 12'b111011101110;
20'b00101001010010101000: color_data = 12'b111011101110;
20'b00101001010010101001: color_data = 12'b111011101110;
20'b00101001010010101010: color_data = 12'b111011101110;
20'b00101001010011101110: color_data = 12'b111011101110;
20'b00101001010011101111: color_data = 12'b111011101110;
20'b00101001010011110000: color_data = 12'b111011101110;
20'b00101001010011110001: color_data = 12'b111011101110;
20'b00101001010011110010: color_data = 12'b111011101110;
20'b00101001010011110011: color_data = 12'b111011101110;
20'b00101001010011110100: color_data = 12'b111011101110;
20'b00101001010011110101: color_data = 12'b111011101110;
20'b00101001010011110110: color_data = 12'b111011101110;
20'b00101001010011110111: color_data = 12'b111011101110;
20'b00101001010011111001: color_data = 12'b111011101110;
20'b00101001010011111010: color_data = 12'b111011101110;
20'b00101001010011111011: color_data = 12'b111011101110;
20'b00101001010011111100: color_data = 12'b111011101110;
20'b00101001010011111101: color_data = 12'b111011101110;
20'b00101001010011111110: color_data = 12'b111011101110;
20'b00101001010011111111: color_data = 12'b111011101110;
20'b00101001010100000000: color_data = 12'b111011101110;
20'b00101001010100000001: color_data = 12'b111011101110;
20'b00101001010100000010: color_data = 12'b111011101110;
20'b00101001010100000100: color_data = 12'b111011101110;
20'b00101001010100000101: color_data = 12'b111011101110;
20'b00101001010100000110: color_data = 12'b111011101110;
20'b00101001010100000111: color_data = 12'b111011101110;
20'b00101001010100001000: color_data = 12'b111011101110;
20'b00101001010100001001: color_data = 12'b111011101110;
20'b00101001010100001010: color_data = 12'b111011101110;
20'b00101001010100001011: color_data = 12'b111011101110;
20'b00101001010100001100: color_data = 12'b111011101110;
20'b00101001010100001101: color_data = 12'b111011101110;
20'b00101001010100001111: color_data = 12'b111011101110;
20'b00101001010100010000: color_data = 12'b111011101110;
20'b00101001010100010001: color_data = 12'b111011101110;
20'b00101001010100010010: color_data = 12'b111011101110;
20'b00101001010100010011: color_data = 12'b111011101110;
20'b00101001010100010100: color_data = 12'b111011101110;
20'b00101001010100010101: color_data = 12'b111011101110;
20'b00101001010100010110: color_data = 12'b111011101110;
20'b00101001010100010111: color_data = 12'b111011101110;
20'b00101001010100011000: color_data = 12'b111011101110;
20'b00101001010100011010: color_data = 12'b111011101110;
20'b00101001010100011011: color_data = 12'b111011101110;
20'b00101001010100011100: color_data = 12'b111011101110;
20'b00101001010100011101: color_data = 12'b111011101110;
20'b00101001010100011110: color_data = 12'b111011101110;
20'b00101001010100011111: color_data = 12'b111011101110;
20'b00101001010100100000: color_data = 12'b111011101110;
20'b00101001010100100001: color_data = 12'b111011101110;
20'b00101001010100100010: color_data = 12'b111011101110;
20'b00101001010100100011: color_data = 12'b111011101110;
20'b00101001010100100101: color_data = 12'b111011101110;
20'b00101001010100100110: color_data = 12'b111011101110;
20'b00101001010100100111: color_data = 12'b111011101110;
20'b00101001010100101000: color_data = 12'b111011101110;
20'b00101001010100101001: color_data = 12'b111011101110;
20'b00101001010100101010: color_data = 12'b111011101110;
20'b00101001010100101011: color_data = 12'b111011101110;
20'b00101001010100101100: color_data = 12'b111011101110;
20'b00101001010100101101: color_data = 12'b111011101110;
20'b00101001010100101110: color_data = 12'b111011101110;
20'b00101001010100110000: color_data = 12'b111011101110;
20'b00101001010100110001: color_data = 12'b111011101110;
20'b00101001010100110010: color_data = 12'b111011101110;
20'b00101001010100110011: color_data = 12'b111011101110;
20'b00101001010100110100: color_data = 12'b111011101110;
20'b00101001010100110101: color_data = 12'b111011101110;
20'b00101001010100110110: color_data = 12'b111011101110;
20'b00101001010100110111: color_data = 12'b111011101110;
20'b00101001010100111000: color_data = 12'b111011101110;
20'b00101001010100111001: color_data = 12'b111011101110;
20'b00101001010101000110: color_data = 12'b111011101110;
20'b00101001010101000111: color_data = 12'b111011101110;
20'b00101001010101001000: color_data = 12'b111011101110;
20'b00101001010101001001: color_data = 12'b111011101110;
20'b00101001010101001010: color_data = 12'b111011101110;
20'b00101001010101001011: color_data = 12'b111011101110;
20'b00101001010101001100: color_data = 12'b111011101110;
20'b00101001010101001101: color_data = 12'b111011101110;
20'b00101001010101001110: color_data = 12'b111011101110;
20'b00101001010101001111: color_data = 12'b111011101110;
20'b00101001010101010001: color_data = 12'b111011101110;
20'b00101001010101010010: color_data = 12'b111011101110;
20'b00101001010101010011: color_data = 12'b111011101110;
20'b00101001010101010100: color_data = 12'b111011101110;
20'b00101001010101010101: color_data = 12'b111011101110;
20'b00101001010101010110: color_data = 12'b111011101110;
20'b00101001010101010111: color_data = 12'b111011101110;
20'b00101001010101011000: color_data = 12'b111011101110;
20'b00101001010101011001: color_data = 12'b111011101110;
20'b00101001010101011010: color_data = 12'b111011101110;
20'b00101001010101111101: color_data = 12'b111011101110;
20'b00101001010101111110: color_data = 12'b111011101110;
20'b00101001010101111111: color_data = 12'b111011101110;
20'b00101001010110000000: color_data = 12'b111011101110;
20'b00101001010110000001: color_data = 12'b111011101110;
20'b00101001010110000010: color_data = 12'b111011101110;
20'b00101001010110000011: color_data = 12'b111011101110;
20'b00101001010110000100: color_data = 12'b111011101110;
20'b00101001010110000101: color_data = 12'b111011101110;
20'b00101001010110000110: color_data = 12'b111011101110;
20'b00101001010110001000: color_data = 12'b111011101110;
20'b00101001010110001001: color_data = 12'b111011101110;
20'b00101001010110001010: color_data = 12'b111011101110;
20'b00101001010110001011: color_data = 12'b111011101110;
20'b00101001010110001100: color_data = 12'b111011101110;
20'b00101001010110001101: color_data = 12'b111011101110;
20'b00101001010110001110: color_data = 12'b111011101110;
20'b00101001010110001111: color_data = 12'b111011101110;
20'b00101001010110010000: color_data = 12'b111011101110;
20'b00101001010110010001: color_data = 12'b111011101110;
20'b00101001010110011110: color_data = 12'b111011101110;
20'b00101001010110011111: color_data = 12'b111011101110;
20'b00101001010110100000: color_data = 12'b111011101110;
20'b00101001010110100001: color_data = 12'b111011101110;
20'b00101001010110100010: color_data = 12'b111011101110;
20'b00101001010110100011: color_data = 12'b111011101110;
20'b00101001010110100100: color_data = 12'b111011101110;
20'b00101001010110100101: color_data = 12'b111011101110;
20'b00101001010110100110: color_data = 12'b111011101110;
20'b00101001010110100111: color_data = 12'b111011101110;
20'b00101001010110101001: color_data = 12'b111011101110;
20'b00101001010110101010: color_data = 12'b111011101110;
20'b00101001010110101011: color_data = 12'b111011101110;
20'b00101001010110101100: color_data = 12'b111011101110;
20'b00101001010110101101: color_data = 12'b111011101110;
20'b00101001010110101110: color_data = 12'b111011101110;
20'b00101001010110101111: color_data = 12'b111011101110;
20'b00101001010110110000: color_data = 12'b111011101110;
20'b00101001010110110001: color_data = 12'b111011101110;
20'b00101001010110110010: color_data = 12'b111011101110;
20'b00101001100011001101: color_data = 12'b111011101110;
20'b00101001100011001110: color_data = 12'b111011101110;
20'b00101001100011001111: color_data = 12'b111011101110;
20'b00101001100011010000: color_data = 12'b111011101110;
20'b00101001100011010001: color_data = 12'b111011101110;
20'b00101001100011010010: color_data = 12'b111011101110;
20'b00101001100011010011: color_data = 12'b111011101110;
20'b00101001100011010100: color_data = 12'b111011101110;
20'b00101001100011010101: color_data = 12'b111011101110;
20'b00101001100011010110: color_data = 12'b111011101110;
20'b00101001100011011000: color_data = 12'b111011101110;
20'b00101001100011011001: color_data = 12'b111011101110;
20'b00101001100011011010: color_data = 12'b111011101110;
20'b00101001100011011011: color_data = 12'b111011101110;
20'b00101001100011011100: color_data = 12'b111011101110;
20'b00101001100011011101: color_data = 12'b111011101110;
20'b00101001100011011110: color_data = 12'b111011101110;
20'b00101001100011011111: color_data = 12'b111011101110;
20'b00101001100011100000: color_data = 12'b111011101110;
20'b00101001100011100001: color_data = 12'b111011101110;
20'b00101001110010010110: color_data = 12'b111011101110;
20'b00101001110010010111: color_data = 12'b111011101110;
20'b00101001110010011000: color_data = 12'b111011101110;
20'b00101001110010011001: color_data = 12'b111011101110;
20'b00101001110010011010: color_data = 12'b111011101110;
20'b00101001110010011011: color_data = 12'b111011101110;
20'b00101001110010011100: color_data = 12'b111011101110;
20'b00101001110010011101: color_data = 12'b111011101110;
20'b00101001110010011110: color_data = 12'b111011101110;
20'b00101001110010011111: color_data = 12'b111011101110;
20'b00101001110010100001: color_data = 12'b111011101110;
20'b00101001110010100010: color_data = 12'b111011101110;
20'b00101001110010100011: color_data = 12'b111011101110;
20'b00101001110010100100: color_data = 12'b111011101110;
20'b00101001110010100101: color_data = 12'b111011101110;
20'b00101001110010100110: color_data = 12'b111011101110;
20'b00101001110010100111: color_data = 12'b111011101110;
20'b00101001110010101000: color_data = 12'b111011101110;
20'b00101001110010101001: color_data = 12'b111011101110;
20'b00101001110010101010: color_data = 12'b111011101110;
20'b00101001110011001101: color_data = 12'b111011101110;
20'b00101001110011001110: color_data = 12'b111011101110;
20'b00101001110011001111: color_data = 12'b111011101110;
20'b00101001110011010000: color_data = 12'b111011101110;
20'b00101001110011010001: color_data = 12'b111011101110;
20'b00101001110011010010: color_data = 12'b111011101110;
20'b00101001110011010011: color_data = 12'b111011101110;
20'b00101001110011010100: color_data = 12'b111011101110;
20'b00101001110011010101: color_data = 12'b111011101110;
20'b00101001110011010110: color_data = 12'b111011101110;
20'b00101001110011011000: color_data = 12'b111011101110;
20'b00101001110011011001: color_data = 12'b111011101110;
20'b00101001110011011010: color_data = 12'b111011101110;
20'b00101001110011011011: color_data = 12'b111011101110;
20'b00101001110011011100: color_data = 12'b111011101110;
20'b00101001110011011101: color_data = 12'b111011101110;
20'b00101001110011011110: color_data = 12'b111011101110;
20'b00101001110011011111: color_data = 12'b111011101110;
20'b00101001110011100000: color_data = 12'b111011101110;
20'b00101001110011100001: color_data = 12'b111011101110;
20'b00101001110011101110: color_data = 12'b111011101110;
20'b00101001110011101111: color_data = 12'b111011101110;
20'b00101001110011110000: color_data = 12'b111011101110;
20'b00101001110011110001: color_data = 12'b111011101110;
20'b00101001110011110010: color_data = 12'b111011101110;
20'b00101001110011110011: color_data = 12'b111011101110;
20'b00101001110011110100: color_data = 12'b111011101110;
20'b00101001110011110101: color_data = 12'b111011101110;
20'b00101001110011110110: color_data = 12'b111011101110;
20'b00101001110011110111: color_data = 12'b111011101110;
20'b00101001110011111001: color_data = 12'b111011101110;
20'b00101001110011111010: color_data = 12'b111011101110;
20'b00101001110011111011: color_data = 12'b111011101110;
20'b00101001110011111100: color_data = 12'b111011101110;
20'b00101001110011111101: color_data = 12'b111011101110;
20'b00101001110011111110: color_data = 12'b111011101110;
20'b00101001110011111111: color_data = 12'b111011101110;
20'b00101001110100000000: color_data = 12'b111011101110;
20'b00101001110100000001: color_data = 12'b111011101110;
20'b00101001110100000010: color_data = 12'b111011101110;
20'b00101001110100100101: color_data = 12'b111011101110;
20'b00101001110100100110: color_data = 12'b111011101110;
20'b00101001110100100111: color_data = 12'b111011101110;
20'b00101001110100101000: color_data = 12'b111011101110;
20'b00101001110100101001: color_data = 12'b111011101110;
20'b00101001110100101010: color_data = 12'b111011101110;
20'b00101001110100101011: color_data = 12'b111011101110;
20'b00101001110100101100: color_data = 12'b111011101110;
20'b00101001110100101101: color_data = 12'b111011101110;
20'b00101001110100101110: color_data = 12'b111011101110;
20'b00101001110100110000: color_data = 12'b111011101110;
20'b00101001110100110001: color_data = 12'b111011101110;
20'b00101001110100110010: color_data = 12'b111011101110;
20'b00101001110100110011: color_data = 12'b111011101110;
20'b00101001110100110100: color_data = 12'b111011101110;
20'b00101001110100110101: color_data = 12'b111011101110;
20'b00101001110100110110: color_data = 12'b111011101110;
20'b00101001110100110111: color_data = 12'b111011101110;
20'b00101001110100111000: color_data = 12'b111011101110;
20'b00101001110100111001: color_data = 12'b111011101110;
20'b00101001110101000110: color_data = 12'b111011101110;
20'b00101001110101000111: color_data = 12'b111011101110;
20'b00101001110101001000: color_data = 12'b111011101110;
20'b00101001110101001001: color_data = 12'b111011101110;
20'b00101001110101001010: color_data = 12'b111011101110;
20'b00101001110101001011: color_data = 12'b111011101110;
20'b00101001110101001100: color_data = 12'b111011101110;
20'b00101001110101001101: color_data = 12'b111011101110;
20'b00101001110101001110: color_data = 12'b111011101110;
20'b00101001110101001111: color_data = 12'b111011101110;
20'b00101001110101010001: color_data = 12'b111011101110;
20'b00101001110101010010: color_data = 12'b111011101110;
20'b00101001110101010011: color_data = 12'b111011101110;
20'b00101001110101010100: color_data = 12'b111011101110;
20'b00101001110101010101: color_data = 12'b111011101110;
20'b00101001110101010110: color_data = 12'b111011101110;
20'b00101001110101010111: color_data = 12'b111011101110;
20'b00101001110101011000: color_data = 12'b111011101110;
20'b00101001110101011001: color_data = 12'b111011101110;
20'b00101001110101011010: color_data = 12'b111011101110;
20'b00101001110101111101: color_data = 12'b111011101110;
20'b00101001110101111110: color_data = 12'b111011101110;
20'b00101001110101111111: color_data = 12'b111011101110;
20'b00101001110110000000: color_data = 12'b111011101110;
20'b00101001110110000001: color_data = 12'b111011101110;
20'b00101001110110000010: color_data = 12'b111011101110;
20'b00101001110110000011: color_data = 12'b111011101110;
20'b00101001110110000100: color_data = 12'b111011101110;
20'b00101001110110000101: color_data = 12'b111011101110;
20'b00101001110110000110: color_data = 12'b111011101110;
20'b00101001110110001000: color_data = 12'b111011101110;
20'b00101001110110001001: color_data = 12'b111011101110;
20'b00101001110110001010: color_data = 12'b111011101110;
20'b00101001110110001011: color_data = 12'b111011101110;
20'b00101001110110001100: color_data = 12'b111011101110;
20'b00101001110110001101: color_data = 12'b111011101110;
20'b00101001110110001110: color_data = 12'b111011101110;
20'b00101001110110001111: color_data = 12'b111011101110;
20'b00101001110110010000: color_data = 12'b111011101110;
20'b00101001110110010001: color_data = 12'b111011101110;
20'b00101001110110011110: color_data = 12'b111011101110;
20'b00101001110110011111: color_data = 12'b111011101110;
20'b00101001110110100000: color_data = 12'b111011101110;
20'b00101001110110100001: color_data = 12'b111011101110;
20'b00101001110110100010: color_data = 12'b111011101110;
20'b00101001110110100011: color_data = 12'b111011101110;
20'b00101001110110100100: color_data = 12'b111011101110;
20'b00101001110110100101: color_data = 12'b111011101110;
20'b00101001110110100110: color_data = 12'b111011101110;
20'b00101001110110100111: color_data = 12'b111011101110;
20'b00101001110110101001: color_data = 12'b111011101110;
20'b00101001110110101010: color_data = 12'b111011101110;
20'b00101001110110101011: color_data = 12'b111011101110;
20'b00101001110110101100: color_data = 12'b111011101110;
20'b00101001110110101101: color_data = 12'b111011101110;
20'b00101001110110101110: color_data = 12'b111011101110;
20'b00101001110110101111: color_data = 12'b111011101110;
20'b00101001110110110000: color_data = 12'b111011101110;
20'b00101001110110110001: color_data = 12'b111011101110;
20'b00101001110110110010: color_data = 12'b111011101110;
20'b00101010000010010110: color_data = 12'b111011101110;
20'b00101010000010010111: color_data = 12'b111011101110;
20'b00101010000010011000: color_data = 12'b111011101110;
20'b00101010000010011001: color_data = 12'b111011101110;
20'b00101010000010011010: color_data = 12'b111011101110;
20'b00101010000010011011: color_data = 12'b111011101110;
20'b00101010000010011100: color_data = 12'b111011101110;
20'b00101010000010011101: color_data = 12'b111011101110;
20'b00101010000010011110: color_data = 12'b111011101110;
20'b00101010000010011111: color_data = 12'b111011101110;
20'b00101010000010100001: color_data = 12'b111011101110;
20'b00101010000010100010: color_data = 12'b111011101110;
20'b00101010000010100011: color_data = 12'b111011101110;
20'b00101010000010100100: color_data = 12'b111011101110;
20'b00101010000010100101: color_data = 12'b111011101110;
20'b00101010000010100110: color_data = 12'b111011101110;
20'b00101010000010100111: color_data = 12'b111011101110;
20'b00101010000010101000: color_data = 12'b111011101110;
20'b00101010000010101001: color_data = 12'b111011101110;
20'b00101010000010101010: color_data = 12'b111011101110;
20'b00101010000011001101: color_data = 12'b111011101110;
20'b00101010000011001110: color_data = 12'b111011101110;
20'b00101010000011001111: color_data = 12'b111011101110;
20'b00101010000011010000: color_data = 12'b111011101110;
20'b00101010000011010001: color_data = 12'b111011101110;
20'b00101010000011010010: color_data = 12'b111011101110;
20'b00101010000011010011: color_data = 12'b111011101110;
20'b00101010000011010100: color_data = 12'b111011101110;
20'b00101010000011010101: color_data = 12'b111011101110;
20'b00101010000011010110: color_data = 12'b111011101110;
20'b00101010000011011000: color_data = 12'b111011101110;
20'b00101010000011011001: color_data = 12'b111011101110;
20'b00101010000011011010: color_data = 12'b111011101110;
20'b00101010000011011011: color_data = 12'b111011101110;
20'b00101010000011011100: color_data = 12'b111011101110;
20'b00101010000011011101: color_data = 12'b111011101110;
20'b00101010000011011110: color_data = 12'b111011101110;
20'b00101010000011011111: color_data = 12'b111011101110;
20'b00101010000011100000: color_data = 12'b111011101110;
20'b00101010000011100001: color_data = 12'b111011101110;
20'b00101010000011101110: color_data = 12'b111011101110;
20'b00101010000011101111: color_data = 12'b111011101110;
20'b00101010000011110000: color_data = 12'b111011101110;
20'b00101010000011110001: color_data = 12'b111011101110;
20'b00101010000011110010: color_data = 12'b111011101110;
20'b00101010000011110011: color_data = 12'b111011101110;
20'b00101010000011110100: color_data = 12'b111011101110;
20'b00101010000011110101: color_data = 12'b111011101110;
20'b00101010000011110110: color_data = 12'b111011101110;
20'b00101010000011110111: color_data = 12'b111011101110;
20'b00101010000011111001: color_data = 12'b111011101110;
20'b00101010000011111010: color_data = 12'b111011101110;
20'b00101010000011111011: color_data = 12'b111011101110;
20'b00101010000011111100: color_data = 12'b111011101110;
20'b00101010000011111101: color_data = 12'b111011101110;
20'b00101010000011111110: color_data = 12'b111011101110;
20'b00101010000011111111: color_data = 12'b111011101110;
20'b00101010000100000000: color_data = 12'b111011101110;
20'b00101010000100000001: color_data = 12'b111011101110;
20'b00101010000100000010: color_data = 12'b111011101110;
20'b00101010000100100101: color_data = 12'b111011101110;
20'b00101010000100100110: color_data = 12'b111011101110;
20'b00101010000100100111: color_data = 12'b111011101110;
20'b00101010000100101000: color_data = 12'b111011101110;
20'b00101010000100101001: color_data = 12'b111011101110;
20'b00101010000100101010: color_data = 12'b111011101110;
20'b00101010000100101011: color_data = 12'b111011101110;
20'b00101010000100101100: color_data = 12'b111011101110;
20'b00101010000100101101: color_data = 12'b111011101110;
20'b00101010000100101110: color_data = 12'b111011101110;
20'b00101010000100110000: color_data = 12'b111011101110;
20'b00101010000100110001: color_data = 12'b111011101110;
20'b00101010000100110010: color_data = 12'b111011101110;
20'b00101010000100110011: color_data = 12'b111011101110;
20'b00101010000100110100: color_data = 12'b111011101110;
20'b00101010000100110101: color_data = 12'b111011101110;
20'b00101010000100110110: color_data = 12'b111011101110;
20'b00101010000100110111: color_data = 12'b111011101110;
20'b00101010000100111000: color_data = 12'b111011101110;
20'b00101010000100111001: color_data = 12'b111011101110;
20'b00101010000101000110: color_data = 12'b111011101110;
20'b00101010000101000111: color_data = 12'b111011101110;
20'b00101010000101001000: color_data = 12'b111011101110;
20'b00101010000101001001: color_data = 12'b111011101110;
20'b00101010000101001010: color_data = 12'b111011101110;
20'b00101010000101001011: color_data = 12'b111011101110;
20'b00101010000101001100: color_data = 12'b111011101110;
20'b00101010000101001101: color_data = 12'b111011101110;
20'b00101010000101001110: color_data = 12'b111011101110;
20'b00101010000101001111: color_data = 12'b111011101110;
20'b00101010000101010001: color_data = 12'b111011101110;
20'b00101010000101010010: color_data = 12'b111011101110;
20'b00101010000101010011: color_data = 12'b111011101110;
20'b00101010000101010100: color_data = 12'b111011101110;
20'b00101010000101010101: color_data = 12'b111011101110;
20'b00101010000101010110: color_data = 12'b111011101110;
20'b00101010000101010111: color_data = 12'b111011101110;
20'b00101010000101011000: color_data = 12'b111011101110;
20'b00101010000101011001: color_data = 12'b111011101110;
20'b00101010000101011010: color_data = 12'b111011101110;
20'b00101010000101111101: color_data = 12'b111011101110;
20'b00101010000101111110: color_data = 12'b111011101110;
20'b00101010000101111111: color_data = 12'b111011101110;
20'b00101010000110000000: color_data = 12'b111011101110;
20'b00101010000110000001: color_data = 12'b111011101110;
20'b00101010000110000010: color_data = 12'b111011101110;
20'b00101010000110000011: color_data = 12'b111011101110;
20'b00101010000110000100: color_data = 12'b111011101110;
20'b00101010000110000101: color_data = 12'b111011101110;
20'b00101010000110000110: color_data = 12'b111011101110;
20'b00101010000110001000: color_data = 12'b111011101110;
20'b00101010000110001001: color_data = 12'b111011101110;
20'b00101010000110001010: color_data = 12'b111011101110;
20'b00101010000110001011: color_data = 12'b111011101110;
20'b00101010000110001100: color_data = 12'b111011101110;
20'b00101010000110001101: color_data = 12'b111011101110;
20'b00101010000110001110: color_data = 12'b111011101110;
20'b00101010000110001111: color_data = 12'b111011101110;
20'b00101010000110010000: color_data = 12'b111011101110;
20'b00101010000110010001: color_data = 12'b111011101110;
20'b00101010000110011110: color_data = 12'b111011101110;
20'b00101010000110011111: color_data = 12'b111011101110;
20'b00101010000110100000: color_data = 12'b111011101110;
20'b00101010000110100001: color_data = 12'b111011101110;
20'b00101010000110100010: color_data = 12'b111011101110;
20'b00101010000110100011: color_data = 12'b111011101110;
20'b00101010000110100100: color_data = 12'b111011101110;
20'b00101010000110100101: color_data = 12'b111011101110;
20'b00101010000110100110: color_data = 12'b111011101110;
20'b00101010000110100111: color_data = 12'b111011101110;
20'b00101010000110101001: color_data = 12'b111011101110;
20'b00101010000110101010: color_data = 12'b111011101110;
20'b00101010000110101011: color_data = 12'b111011101110;
20'b00101010000110101100: color_data = 12'b111011101110;
20'b00101010000110101101: color_data = 12'b111011101110;
20'b00101010000110101110: color_data = 12'b111011101110;
20'b00101010000110101111: color_data = 12'b111011101110;
20'b00101010000110110000: color_data = 12'b111011101110;
20'b00101010000110110001: color_data = 12'b111011101110;
20'b00101010000110110010: color_data = 12'b111011101110;
20'b00101010010010010110: color_data = 12'b111011101110;
20'b00101010010010010111: color_data = 12'b111011101110;
20'b00101010010010011000: color_data = 12'b111011101110;
20'b00101010010010011001: color_data = 12'b111011101110;
20'b00101010010010011010: color_data = 12'b111011101110;
20'b00101010010010011011: color_data = 12'b111011101110;
20'b00101010010010011100: color_data = 12'b111011101110;
20'b00101010010010011101: color_data = 12'b111011101110;
20'b00101010010010011110: color_data = 12'b111011101110;
20'b00101010010010011111: color_data = 12'b111011101110;
20'b00101010010010100001: color_data = 12'b111011101110;
20'b00101010010010100010: color_data = 12'b111011101110;
20'b00101010010010100011: color_data = 12'b111011101110;
20'b00101010010010100100: color_data = 12'b111011101110;
20'b00101010010010100101: color_data = 12'b111011101110;
20'b00101010010010100110: color_data = 12'b111011101110;
20'b00101010010010100111: color_data = 12'b111011101110;
20'b00101010010010101000: color_data = 12'b111011101110;
20'b00101010010010101001: color_data = 12'b111011101110;
20'b00101010010010101010: color_data = 12'b111011101110;
20'b00101010010011001101: color_data = 12'b111011101110;
20'b00101010010011001110: color_data = 12'b111011101110;
20'b00101010010011001111: color_data = 12'b111011101110;
20'b00101010010011010000: color_data = 12'b111011101110;
20'b00101010010011010001: color_data = 12'b111011101110;
20'b00101010010011010010: color_data = 12'b111011101110;
20'b00101010010011010011: color_data = 12'b111011101110;
20'b00101010010011010100: color_data = 12'b111011101110;
20'b00101010010011010101: color_data = 12'b111011101110;
20'b00101010010011010110: color_data = 12'b111011101110;
20'b00101010010011011000: color_data = 12'b111011101110;
20'b00101010010011011001: color_data = 12'b111011101110;
20'b00101010010011011010: color_data = 12'b111011101110;
20'b00101010010011011011: color_data = 12'b111011101110;
20'b00101010010011011100: color_data = 12'b111011101110;
20'b00101010010011011101: color_data = 12'b111011101110;
20'b00101010010011011110: color_data = 12'b111011101110;
20'b00101010010011011111: color_data = 12'b111011101110;
20'b00101010010011100000: color_data = 12'b111011101110;
20'b00101010010011100001: color_data = 12'b111011101110;
20'b00101010010011101110: color_data = 12'b111011101110;
20'b00101010010011101111: color_data = 12'b111011101110;
20'b00101010010011110000: color_data = 12'b111011101110;
20'b00101010010011110001: color_data = 12'b111011101110;
20'b00101010010011110010: color_data = 12'b111011101110;
20'b00101010010011110011: color_data = 12'b111011101110;
20'b00101010010011110100: color_data = 12'b111011101110;
20'b00101010010011110101: color_data = 12'b111011101110;
20'b00101010010011110110: color_data = 12'b111011101110;
20'b00101010010011110111: color_data = 12'b111011101110;
20'b00101010010011111001: color_data = 12'b111011101110;
20'b00101010010011111010: color_data = 12'b111011101110;
20'b00101010010011111011: color_data = 12'b111011101110;
20'b00101010010011111100: color_data = 12'b111011101110;
20'b00101010010011111101: color_data = 12'b111011101110;
20'b00101010010011111110: color_data = 12'b111011101110;
20'b00101010010011111111: color_data = 12'b111011101110;
20'b00101010010100000000: color_data = 12'b111011101110;
20'b00101010010100000001: color_data = 12'b111011101110;
20'b00101010010100000010: color_data = 12'b111011101110;
20'b00101010010100100101: color_data = 12'b111011101110;
20'b00101010010100100110: color_data = 12'b111011101110;
20'b00101010010100100111: color_data = 12'b111011101110;
20'b00101010010100101000: color_data = 12'b111011101110;
20'b00101010010100101001: color_data = 12'b111011101110;
20'b00101010010100101010: color_data = 12'b111011101110;
20'b00101010010100101011: color_data = 12'b111011101110;
20'b00101010010100101100: color_data = 12'b111011101110;
20'b00101010010100101101: color_data = 12'b111011101110;
20'b00101010010100101110: color_data = 12'b111011101110;
20'b00101010010100110000: color_data = 12'b111011101110;
20'b00101010010100110001: color_data = 12'b111011101110;
20'b00101010010100110010: color_data = 12'b111011101110;
20'b00101010010100110011: color_data = 12'b111011101110;
20'b00101010010100110100: color_data = 12'b111011101110;
20'b00101010010100110101: color_data = 12'b111011101110;
20'b00101010010100110110: color_data = 12'b111011101110;
20'b00101010010100110111: color_data = 12'b111011101110;
20'b00101010010100111000: color_data = 12'b111011101110;
20'b00101010010100111001: color_data = 12'b111011101110;
20'b00101010010101000110: color_data = 12'b111011101110;
20'b00101010010101000111: color_data = 12'b111011101110;
20'b00101010010101001000: color_data = 12'b111011101110;
20'b00101010010101001001: color_data = 12'b111011101110;
20'b00101010010101001010: color_data = 12'b111011101110;
20'b00101010010101001011: color_data = 12'b111011101110;
20'b00101010010101001100: color_data = 12'b111011101110;
20'b00101010010101001101: color_data = 12'b111011101110;
20'b00101010010101001110: color_data = 12'b111011101110;
20'b00101010010101001111: color_data = 12'b111011101110;
20'b00101010010101010001: color_data = 12'b111011101110;
20'b00101010010101010010: color_data = 12'b111011101110;
20'b00101010010101010011: color_data = 12'b111011101110;
20'b00101010010101010100: color_data = 12'b111011101110;
20'b00101010010101010101: color_data = 12'b111011101110;
20'b00101010010101010110: color_data = 12'b111011101110;
20'b00101010010101010111: color_data = 12'b111011101110;
20'b00101010010101011000: color_data = 12'b111011101110;
20'b00101010010101011001: color_data = 12'b111011101110;
20'b00101010010101011010: color_data = 12'b111011101110;
20'b00101010010101111101: color_data = 12'b111011101110;
20'b00101010010101111110: color_data = 12'b111011101110;
20'b00101010010101111111: color_data = 12'b111011101110;
20'b00101010010110000000: color_data = 12'b111011101110;
20'b00101010010110000001: color_data = 12'b111011101110;
20'b00101010010110000010: color_data = 12'b111011101110;
20'b00101010010110000011: color_data = 12'b111011101110;
20'b00101010010110000100: color_data = 12'b111011101110;
20'b00101010010110000101: color_data = 12'b111011101110;
20'b00101010010110000110: color_data = 12'b111011101110;
20'b00101010010110001000: color_data = 12'b111011101110;
20'b00101010010110001001: color_data = 12'b111011101110;
20'b00101010010110001010: color_data = 12'b111011101110;
20'b00101010010110001011: color_data = 12'b111011101110;
20'b00101010010110001100: color_data = 12'b111011101110;
20'b00101010010110001101: color_data = 12'b111011101110;
20'b00101010010110001110: color_data = 12'b111011101110;
20'b00101010010110001111: color_data = 12'b111011101110;
20'b00101010010110010000: color_data = 12'b111011101110;
20'b00101010010110010001: color_data = 12'b111011101110;
20'b00101010010110011110: color_data = 12'b111011101110;
20'b00101010010110011111: color_data = 12'b111011101110;
20'b00101010010110100000: color_data = 12'b111011101110;
20'b00101010010110100001: color_data = 12'b111011101110;
20'b00101010010110100010: color_data = 12'b111011101110;
20'b00101010010110100011: color_data = 12'b111011101110;
20'b00101010010110100100: color_data = 12'b111011101110;
20'b00101010010110100101: color_data = 12'b111011101110;
20'b00101010010110100110: color_data = 12'b111011101110;
20'b00101010010110100111: color_data = 12'b111011101110;
20'b00101010010110101001: color_data = 12'b111011101110;
20'b00101010010110101010: color_data = 12'b111011101110;
20'b00101010010110101011: color_data = 12'b111011101110;
20'b00101010010110101100: color_data = 12'b111011101110;
20'b00101010010110101101: color_data = 12'b111011101110;
20'b00101010010110101110: color_data = 12'b111011101110;
20'b00101010010110101111: color_data = 12'b111011101110;
20'b00101010010110110000: color_data = 12'b111011101110;
20'b00101010010110110001: color_data = 12'b111011101110;
20'b00101010010110110010: color_data = 12'b111011101110;
20'b00101010100010010110: color_data = 12'b111011101110;
20'b00101010100010010111: color_data = 12'b111011101110;
20'b00101010100010011000: color_data = 12'b111011101110;
20'b00101010100010011001: color_data = 12'b111011101110;
20'b00101010100010011010: color_data = 12'b111011101110;
20'b00101010100010011011: color_data = 12'b111011101110;
20'b00101010100010011100: color_data = 12'b111011101110;
20'b00101010100010011101: color_data = 12'b111011101110;
20'b00101010100010011110: color_data = 12'b111011101110;
20'b00101010100010011111: color_data = 12'b111011101110;
20'b00101010100010100001: color_data = 12'b111011101110;
20'b00101010100010100010: color_data = 12'b111011101110;
20'b00101010100010100011: color_data = 12'b111011101110;
20'b00101010100010100100: color_data = 12'b111011101110;
20'b00101010100010100101: color_data = 12'b111011101110;
20'b00101010100010100110: color_data = 12'b111011101110;
20'b00101010100010100111: color_data = 12'b111011101110;
20'b00101010100010101000: color_data = 12'b111011101110;
20'b00101010100010101001: color_data = 12'b111011101110;
20'b00101010100010101010: color_data = 12'b111011101110;
20'b00101010100011001101: color_data = 12'b111011101110;
20'b00101010100011001110: color_data = 12'b111011101110;
20'b00101010100011001111: color_data = 12'b111011101110;
20'b00101010100011010000: color_data = 12'b111011101110;
20'b00101010100011010001: color_data = 12'b111011101110;
20'b00101010100011010010: color_data = 12'b111011101110;
20'b00101010100011010011: color_data = 12'b111011101110;
20'b00101010100011010100: color_data = 12'b111011101110;
20'b00101010100011010101: color_data = 12'b111011101110;
20'b00101010100011010110: color_data = 12'b111011101110;
20'b00101010100011011000: color_data = 12'b111011101110;
20'b00101010100011011001: color_data = 12'b111011101110;
20'b00101010100011011010: color_data = 12'b111011101110;
20'b00101010100011011011: color_data = 12'b111011101110;
20'b00101010100011011100: color_data = 12'b111011101110;
20'b00101010100011011101: color_data = 12'b111011101110;
20'b00101010100011011110: color_data = 12'b111011101110;
20'b00101010100011011111: color_data = 12'b111011101110;
20'b00101010100011100000: color_data = 12'b111011101110;
20'b00101010100011100001: color_data = 12'b111011101110;
20'b00101010100011101110: color_data = 12'b111011101110;
20'b00101010100011101111: color_data = 12'b111011101110;
20'b00101010100011110000: color_data = 12'b111011101110;
20'b00101010100011110001: color_data = 12'b111011101110;
20'b00101010100011110010: color_data = 12'b111011101110;
20'b00101010100011110011: color_data = 12'b111011101110;
20'b00101010100011110100: color_data = 12'b111011101110;
20'b00101010100011110101: color_data = 12'b111011101110;
20'b00101010100011110110: color_data = 12'b111011101110;
20'b00101010100011110111: color_data = 12'b111011101110;
20'b00101010100011111001: color_data = 12'b111011101110;
20'b00101010100011111010: color_data = 12'b111011101110;
20'b00101010100011111011: color_data = 12'b111011101110;
20'b00101010100011111100: color_data = 12'b111011101110;
20'b00101010100011111101: color_data = 12'b111011101110;
20'b00101010100011111110: color_data = 12'b111011101110;
20'b00101010100011111111: color_data = 12'b111011101110;
20'b00101010100100000000: color_data = 12'b111011101110;
20'b00101010100100000001: color_data = 12'b111011101110;
20'b00101010100100000010: color_data = 12'b111011101110;
20'b00101010100100100101: color_data = 12'b111011101110;
20'b00101010100100100110: color_data = 12'b111011101110;
20'b00101010100100100111: color_data = 12'b111011101110;
20'b00101010100100101000: color_data = 12'b111011101110;
20'b00101010100100101001: color_data = 12'b111011101110;
20'b00101010100100101010: color_data = 12'b111011101110;
20'b00101010100100101011: color_data = 12'b111011101110;
20'b00101010100100101100: color_data = 12'b111011101110;
20'b00101010100100101101: color_data = 12'b111011101110;
20'b00101010100100101110: color_data = 12'b111011101110;
20'b00101010100100110000: color_data = 12'b111011101110;
20'b00101010100100110001: color_data = 12'b111011101110;
20'b00101010100100110010: color_data = 12'b111011101110;
20'b00101010100100110011: color_data = 12'b111011101110;
20'b00101010100100110100: color_data = 12'b111011101110;
20'b00101010100100110101: color_data = 12'b111011101110;
20'b00101010100100110110: color_data = 12'b111011101110;
20'b00101010100100110111: color_data = 12'b111011101110;
20'b00101010100100111000: color_data = 12'b111011101110;
20'b00101010100100111001: color_data = 12'b111011101110;
20'b00101010100101000110: color_data = 12'b111011101110;
20'b00101010100101000111: color_data = 12'b111011101110;
20'b00101010100101001000: color_data = 12'b111011101110;
20'b00101010100101001001: color_data = 12'b111011101110;
20'b00101010100101001010: color_data = 12'b111011101110;
20'b00101010100101001011: color_data = 12'b111011101110;
20'b00101010100101001100: color_data = 12'b111011101110;
20'b00101010100101001101: color_data = 12'b111011101110;
20'b00101010100101001110: color_data = 12'b111011101110;
20'b00101010100101001111: color_data = 12'b111011101110;
20'b00101010100101010001: color_data = 12'b111011101110;
20'b00101010100101010010: color_data = 12'b111011101110;
20'b00101010100101010011: color_data = 12'b111011101110;
20'b00101010100101010100: color_data = 12'b111011101110;
20'b00101010100101010101: color_data = 12'b111011101110;
20'b00101010100101010110: color_data = 12'b111011101110;
20'b00101010100101010111: color_data = 12'b111011101110;
20'b00101010100101011000: color_data = 12'b111011101110;
20'b00101010100101011001: color_data = 12'b111011101110;
20'b00101010100101011010: color_data = 12'b111011101110;
20'b00101010100101111101: color_data = 12'b111011101110;
20'b00101010100101111110: color_data = 12'b111011101110;
20'b00101010100101111111: color_data = 12'b111011101110;
20'b00101010100110000000: color_data = 12'b111011101110;
20'b00101010100110000001: color_data = 12'b111011101110;
20'b00101010100110000010: color_data = 12'b111011101110;
20'b00101010100110000011: color_data = 12'b111011101110;
20'b00101010100110000100: color_data = 12'b111011101110;
20'b00101010100110000101: color_data = 12'b111011101110;
20'b00101010100110000110: color_data = 12'b111011101110;
20'b00101010100110001000: color_data = 12'b111011101110;
20'b00101010100110001001: color_data = 12'b111011101110;
20'b00101010100110001010: color_data = 12'b111011101110;
20'b00101010100110001011: color_data = 12'b111011101110;
20'b00101010100110001100: color_data = 12'b111011101110;
20'b00101010100110001101: color_data = 12'b111011101110;
20'b00101010100110001110: color_data = 12'b111011101110;
20'b00101010100110001111: color_data = 12'b111011101110;
20'b00101010100110010000: color_data = 12'b111011101110;
20'b00101010100110010001: color_data = 12'b111011101110;
20'b00101010100110011110: color_data = 12'b111011101110;
20'b00101010100110011111: color_data = 12'b111011101110;
20'b00101010100110100000: color_data = 12'b111011101110;
20'b00101010100110100001: color_data = 12'b111011101110;
20'b00101010100110100010: color_data = 12'b111011101110;
20'b00101010100110100011: color_data = 12'b111011101110;
20'b00101010100110100100: color_data = 12'b111011101110;
20'b00101010100110100101: color_data = 12'b111011101110;
20'b00101010100110100110: color_data = 12'b111011101110;
20'b00101010100110100111: color_data = 12'b111011101110;
20'b00101010100110101001: color_data = 12'b111011101110;
20'b00101010100110101010: color_data = 12'b111011101110;
20'b00101010100110101011: color_data = 12'b111011101110;
20'b00101010100110101100: color_data = 12'b111011101110;
20'b00101010100110101101: color_data = 12'b111011101110;
20'b00101010100110101110: color_data = 12'b111011101110;
20'b00101010100110101111: color_data = 12'b111011101110;
20'b00101010100110110000: color_data = 12'b111011101110;
20'b00101010100110110001: color_data = 12'b111011101110;
20'b00101010100110110010: color_data = 12'b111011101110;
20'b00101010110010010110: color_data = 12'b111011101110;
20'b00101010110010010111: color_data = 12'b111011101110;
20'b00101010110010011000: color_data = 12'b111011101110;
20'b00101010110010011001: color_data = 12'b111011101110;
20'b00101010110010011010: color_data = 12'b111011101110;
20'b00101010110010011011: color_data = 12'b111011101110;
20'b00101010110010011100: color_data = 12'b111011101110;
20'b00101010110010011101: color_data = 12'b111011101110;
20'b00101010110010011110: color_data = 12'b111011101110;
20'b00101010110010011111: color_data = 12'b111011101110;
20'b00101010110010100001: color_data = 12'b111011101110;
20'b00101010110010100010: color_data = 12'b111011101110;
20'b00101010110010100011: color_data = 12'b111011101110;
20'b00101010110010100100: color_data = 12'b111011101110;
20'b00101010110010100101: color_data = 12'b111011101110;
20'b00101010110010100110: color_data = 12'b111011101110;
20'b00101010110010100111: color_data = 12'b111011101110;
20'b00101010110010101000: color_data = 12'b111011101110;
20'b00101010110010101001: color_data = 12'b111011101110;
20'b00101010110010101010: color_data = 12'b111011101110;
20'b00101010110011001101: color_data = 12'b111011101110;
20'b00101010110011001110: color_data = 12'b111011101110;
20'b00101010110011001111: color_data = 12'b111011101110;
20'b00101010110011010000: color_data = 12'b111011101110;
20'b00101010110011010001: color_data = 12'b111011101110;
20'b00101010110011010010: color_data = 12'b111011101110;
20'b00101010110011010011: color_data = 12'b111011101110;
20'b00101010110011010100: color_data = 12'b111011101110;
20'b00101010110011010101: color_data = 12'b111011101110;
20'b00101010110011010110: color_data = 12'b111011101110;
20'b00101010110011011000: color_data = 12'b111011101110;
20'b00101010110011011001: color_data = 12'b111011101110;
20'b00101010110011011010: color_data = 12'b111011101110;
20'b00101010110011011011: color_data = 12'b111011101110;
20'b00101010110011011100: color_data = 12'b111011101110;
20'b00101010110011011101: color_data = 12'b111011101110;
20'b00101010110011011110: color_data = 12'b111011101110;
20'b00101010110011011111: color_data = 12'b111011101110;
20'b00101010110011100000: color_data = 12'b111011101110;
20'b00101010110011100001: color_data = 12'b111011101110;
20'b00101010110011101110: color_data = 12'b111011101110;
20'b00101010110011101111: color_data = 12'b111011101110;
20'b00101010110011110000: color_data = 12'b111011101110;
20'b00101010110011110001: color_data = 12'b111011101110;
20'b00101010110011110010: color_data = 12'b111011101110;
20'b00101010110011110011: color_data = 12'b111011101110;
20'b00101010110011110100: color_data = 12'b111011101110;
20'b00101010110011110101: color_data = 12'b111011101110;
20'b00101010110011110110: color_data = 12'b111011101110;
20'b00101010110011110111: color_data = 12'b111011101110;
20'b00101010110011111001: color_data = 12'b111011101110;
20'b00101010110011111010: color_data = 12'b111011101110;
20'b00101010110011111011: color_data = 12'b111011101110;
20'b00101010110011111100: color_data = 12'b111011101110;
20'b00101010110011111101: color_data = 12'b111011101110;
20'b00101010110011111110: color_data = 12'b111011101110;
20'b00101010110011111111: color_data = 12'b111011101110;
20'b00101010110100000000: color_data = 12'b111011101110;
20'b00101010110100000001: color_data = 12'b111011101110;
20'b00101010110100000010: color_data = 12'b111011101110;
20'b00101010110100100101: color_data = 12'b111011101110;
20'b00101010110100100110: color_data = 12'b111011101110;
20'b00101010110100100111: color_data = 12'b111011101110;
20'b00101010110100101000: color_data = 12'b111011101110;
20'b00101010110100101001: color_data = 12'b111011101110;
20'b00101010110100101010: color_data = 12'b111011101110;
20'b00101010110100101011: color_data = 12'b111011101110;
20'b00101010110100101100: color_data = 12'b111011101110;
20'b00101010110100101101: color_data = 12'b111011101110;
20'b00101010110100101110: color_data = 12'b111011101110;
20'b00101010110100110000: color_data = 12'b111011101110;
20'b00101010110100110001: color_data = 12'b111011101110;
20'b00101010110100110010: color_data = 12'b111011101110;
20'b00101010110100110011: color_data = 12'b111011101110;
20'b00101010110100110100: color_data = 12'b111011101110;
20'b00101010110100110101: color_data = 12'b111011101110;
20'b00101010110100110110: color_data = 12'b111011101110;
20'b00101010110100110111: color_data = 12'b111011101110;
20'b00101010110100111000: color_data = 12'b111011101110;
20'b00101010110100111001: color_data = 12'b111011101110;
20'b00101010110101000110: color_data = 12'b111011101110;
20'b00101010110101000111: color_data = 12'b111011101110;
20'b00101010110101001000: color_data = 12'b111011101110;
20'b00101010110101001001: color_data = 12'b111011101110;
20'b00101010110101001010: color_data = 12'b111011101110;
20'b00101010110101001011: color_data = 12'b111011101110;
20'b00101010110101001100: color_data = 12'b111011101110;
20'b00101010110101001101: color_data = 12'b111011101110;
20'b00101010110101001110: color_data = 12'b111011101110;
20'b00101010110101001111: color_data = 12'b111011101110;
20'b00101010110101010001: color_data = 12'b111011101110;
20'b00101010110101010010: color_data = 12'b111011101110;
20'b00101010110101010011: color_data = 12'b111011101110;
20'b00101010110101010100: color_data = 12'b111011101110;
20'b00101010110101010101: color_data = 12'b111011101110;
20'b00101010110101010110: color_data = 12'b111011101110;
20'b00101010110101010111: color_data = 12'b111011101110;
20'b00101010110101011000: color_data = 12'b111011101110;
20'b00101010110101011001: color_data = 12'b111011101110;
20'b00101010110101011010: color_data = 12'b111011101110;
20'b00101010110101111101: color_data = 12'b111011101110;
20'b00101010110101111110: color_data = 12'b111011101110;
20'b00101010110101111111: color_data = 12'b111011101110;
20'b00101010110110000000: color_data = 12'b111011101110;
20'b00101010110110000001: color_data = 12'b111011101110;
20'b00101010110110000010: color_data = 12'b111011101110;
20'b00101010110110000011: color_data = 12'b111011101110;
20'b00101010110110000100: color_data = 12'b111011101110;
20'b00101010110110000101: color_data = 12'b111011101110;
20'b00101010110110000110: color_data = 12'b111011101110;
20'b00101010110110001000: color_data = 12'b111011101110;
20'b00101010110110001001: color_data = 12'b111011101110;
20'b00101010110110001010: color_data = 12'b111011101110;
20'b00101010110110001011: color_data = 12'b111011101110;
20'b00101010110110001100: color_data = 12'b111011101110;
20'b00101010110110001101: color_data = 12'b111011101110;
20'b00101010110110001110: color_data = 12'b111011101110;
20'b00101010110110001111: color_data = 12'b111011101110;
20'b00101010110110010000: color_data = 12'b111011101110;
20'b00101010110110010001: color_data = 12'b111011101110;
20'b00101010110110011110: color_data = 12'b111011101110;
20'b00101010110110011111: color_data = 12'b111011101110;
20'b00101010110110100000: color_data = 12'b111011101110;
20'b00101010110110100001: color_data = 12'b111011101110;
20'b00101010110110100010: color_data = 12'b111011101110;
20'b00101010110110100011: color_data = 12'b111011101110;
20'b00101010110110100100: color_data = 12'b111011101110;
20'b00101010110110100101: color_data = 12'b111011101110;
20'b00101010110110100110: color_data = 12'b111011101110;
20'b00101010110110100111: color_data = 12'b111011101110;
20'b00101010110110101001: color_data = 12'b111011101110;
20'b00101010110110101010: color_data = 12'b111011101110;
20'b00101010110110101011: color_data = 12'b111011101110;
20'b00101010110110101100: color_data = 12'b111011101110;
20'b00101010110110101101: color_data = 12'b111011101110;
20'b00101010110110101110: color_data = 12'b111011101110;
20'b00101010110110101111: color_data = 12'b111011101110;
20'b00101010110110110000: color_data = 12'b111011101110;
20'b00101010110110110001: color_data = 12'b111011101110;
20'b00101010110110110010: color_data = 12'b111011101110;
20'b00101011000010010110: color_data = 12'b111011101110;
20'b00101011000010010111: color_data = 12'b111011101110;
20'b00101011000010011000: color_data = 12'b111011101110;
20'b00101011000010011001: color_data = 12'b111011101110;
20'b00101011000010011010: color_data = 12'b111011101110;
20'b00101011000010011011: color_data = 12'b111011101110;
20'b00101011000010011100: color_data = 12'b111011101110;
20'b00101011000010011101: color_data = 12'b111011101110;
20'b00101011000010011110: color_data = 12'b111011101110;
20'b00101011000010011111: color_data = 12'b111011101110;
20'b00101011000010100001: color_data = 12'b111011101110;
20'b00101011000010100010: color_data = 12'b111011101110;
20'b00101011000010100011: color_data = 12'b111011101110;
20'b00101011000010100100: color_data = 12'b111011101110;
20'b00101011000010100101: color_data = 12'b111011101110;
20'b00101011000010100110: color_data = 12'b111011101110;
20'b00101011000010100111: color_data = 12'b111011101110;
20'b00101011000010101000: color_data = 12'b111011101110;
20'b00101011000010101001: color_data = 12'b111011101110;
20'b00101011000010101010: color_data = 12'b111011101110;
20'b00101011000011001101: color_data = 12'b111011101110;
20'b00101011000011001110: color_data = 12'b111011101110;
20'b00101011000011001111: color_data = 12'b111011101110;
20'b00101011000011010000: color_data = 12'b111011101110;
20'b00101011000011010001: color_data = 12'b111011101110;
20'b00101011000011010010: color_data = 12'b111011101110;
20'b00101011000011010011: color_data = 12'b111011101110;
20'b00101011000011010100: color_data = 12'b111011101110;
20'b00101011000011010101: color_data = 12'b111011101110;
20'b00101011000011010110: color_data = 12'b111011101110;
20'b00101011000011011000: color_data = 12'b111011101110;
20'b00101011000011011001: color_data = 12'b111011101110;
20'b00101011000011011010: color_data = 12'b111011101110;
20'b00101011000011011011: color_data = 12'b111011101110;
20'b00101011000011011100: color_data = 12'b111011101110;
20'b00101011000011011101: color_data = 12'b111011101110;
20'b00101011000011011110: color_data = 12'b111011101110;
20'b00101011000011011111: color_data = 12'b111011101110;
20'b00101011000011100000: color_data = 12'b111011101110;
20'b00101011000011100001: color_data = 12'b111011101110;
20'b00101011000011101110: color_data = 12'b111011101110;
20'b00101011000011101111: color_data = 12'b111011101110;
20'b00101011000011110000: color_data = 12'b111011101110;
20'b00101011000011110001: color_data = 12'b111011101110;
20'b00101011000011110010: color_data = 12'b111011101110;
20'b00101011000011110011: color_data = 12'b111011101110;
20'b00101011000011110100: color_data = 12'b111011101110;
20'b00101011000011110101: color_data = 12'b111011101110;
20'b00101011000011110110: color_data = 12'b111011101110;
20'b00101011000011110111: color_data = 12'b111011101110;
20'b00101011000011111001: color_data = 12'b111011101110;
20'b00101011000011111010: color_data = 12'b111011101110;
20'b00101011000011111011: color_data = 12'b111011101110;
20'b00101011000011111100: color_data = 12'b111011101110;
20'b00101011000011111101: color_data = 12'b111011101110;
20'b00101011000011111110: color_data = 12'b111011101110;
20'b00101011000011111111: color_data = 12'b111011101110;
20'b00101011000100000000: color_data = 12'b111011101110;
20'b00101011000100000001: color_data = 12'b111011101110;
20'b00101011000100000010: color_data = 12'b111011101110;
20'b00101011000100100101: color_data = 12'b111011101110;
20'b00101011000100100110: color_data = 12'b111011101110;
20'b00101011000100100111: color_data = 12'b111011101110;
20'b00101011000100101000: color_data = 12'b111011101110;
20'b00101011000100101001: color_data = 12'b111011101110;
20'b00101011000100101010: color_data = 12'b111011101110;
20'b00101011000100101011: color_data = 12'b111011101110;
20'b00101011000100101100: color_data = 12'b111011101110;
20'b00101011000100101101: color_data = 12'b111011101110;
20'b00101011000100101110: color_data = 12'b111011101110;
20'b00101011000100110000: color_data = 12'b111011101110;
20'b00101011000100110001: color_data = 12'b111011101110;
20'b00101011000100110010: color_data = 12'b111011101110;
20'b00101011000100110011: color_data = 12'b111011101110;
20'b00101011000100110100: color_data = 12'b111011101110;
20'b00101011000100110101: color_data = 12'b111011101110;
20'b00101011000100110110: color_data = 12'b111011101110;
20'b00101011000100110111: color_data = 12'b111011101110;
20'b00101011000100111000: color_data = 12'b111011101110;
20'b00101011000100111001: color_data = 12'b111011101110;
20'b00101011000101000110: color_data = 12'b111011101110;
20'b00101011000101000111: color_data = 12'b111011101110;
20'b00101011000101001000: color_data = 12'b111011101110;
20'b00101011000101001001: color_data = 12'b111011101110;
20'b00101011000101001010: color_data = 12'b111011101110;
20'b00101011000101001011: color_data = 12'b111011101110;
20'b00101011000101001100: color_data = 12'b111011101110;
20'b00101011000101001101: color_data = 12'b111011101110;
20'b00101011000101001110: color_data = 12'b111011101110;
20'b00101011000101001111: color_data = 12'b111011101110;
20'b00101011000101010001: color_data = 12'b111011101110;
20'b00101011000101010010: color_data = 12'b111011101110;
20'b00101011000101010011: color_data = 12'b111011101110;
20'b00101011000101010100: color_data = 12'b111011101110;
20'b00101011000101010101: color_data = 12'b111011101110;
20'b00101011000101010110: color_data = 12'b111011101110;
20'b00101011000101010111: color_data = 12'b111011101110;
20'b00101011000101011000: color_data = 12'b111011101110;
20'b00101011000101011001: color_data = 12'b111011101110;
20'b00101011000101011010: color_data = 12'b111011101110;
20'b00101011000101111101: color_data = 12'b111011101110;
20'b00101011000101111110: color_data = 12'b111011101110;
20'b00101011000101111111: color_data = 12'b111011101110;
20'b00101011000110000000: color_data = 12'b111011101110;
20'b00101011000110000001: color_data = 12'b111011101110;
20'b00101011000110000010: color_data = 12'b111011101110;
20'b00101011000110000011: color_data = 12'b111011101110;
20'b00101011000110000100: color_data = 12'b111011101110;
20'b00101011000110000101: color_data = 12'b111011101110;
20'b00101011000110000110: color_data = 12'b111011101110;
20'b00101011000110001000: color_data = 12'b111011101110;
20'b00101011000110001001: color_data = 12'b111011101110;
20'b00101011000110001010: color_data = 12'b111011101110;
20'b00101011000110001011: color_data = 12'b111011101110;
20'b00101011000110001100: color_data = 12'b111011101110;
20'b00101011000110001101: color_data = 12'b111011101110;
20'b00101011000110001110: color_data = 12'b111011101110;
20'b00101011000110001111: color_data = 12'b111011101110;
20'b00101011000110010000: color_data = 12'b111011101110;
20'b00101011000110010001: color_data = 12'b111011101110;
20'b00101011000110011110: color_data = 12'b111011101110;
20'b00101011000110011111: color_data = 12'b111011101110;
20'b00101011000110100000: color_data = 12'b111011101110;
20'b00101011000110100001: color_data = 12'b111011101110;
20'b00101011000110100010: color_data = 12'b111011101110;
20'b00101011000110100011: color_data = 12'b111011101110;
20'b00101011000110100100: color_data = 12'b111011101110;
20'b00101011000110100101: color_data = 12'b111011101110;
20'b00101011000110100110: color_data = 12'b111011101110;
20'b00101011000110100111: color_data = 12'b111011101110;
20'b00101011000110101001: color_data = 12'b111011101110;
20'b00101011000110101010: color_data = 12'b111011101110;
20'b00101011000110101011: color_data = 12'b111011101110;
20'b00101011000110101100: color_data = 12'b111011101110;
20'b00101011000110101101: color_data = 12'b111011101110;
20'b00101011000110101110: color_data = 12'b111011101110;
20'b00101011000110101111: color_data = 12'b111011101110;
20'b00101011000110110000: color_data = 12'b111011101110;
20'b00101011000110110001: color_data = 12'b111011101110;
20'b00101011000110110010: color_data = 12'b111011101110;
20'b00101011010010010110: color_data = 12'b111011101110;
20'b00101011010010010111: color_data = 12'b111011101110;
20'b00101011010010011000: color_data = 12'b111011101110;
20'b00101011010010011001: color_data = 12'b111011101110;
20'b00101011010010011010: color_data = 12'b111011101110;
20'b00101011010010011011: color_data = 12'b111011101110;
20'b00101011010010011100: color_data = 12'b111011101110;
20'b00101011010010011101: color_data = 12'b111011101110;
20'b00101011010010011110: color_data = 12'b111011101110;
20'b00101011010010011111: color_data = 12'b111011101110;
20'b00101011010010100001: color_data = 12'b111011101110;
20'b00101011010010100010: color_data = 12'b111011101110;
20'b00101011010010100011: color_data = 12'b111011101110;
20'b00101011010010100100: color_data = 12'b111011101110;
20'b00101011010010100101: color_data = 12'b111011101110;
20'b00101011010010100110: color_data = 12'b111011101110;
20'b00101011010010100111: color_data = 12'b111011101110;
20'b00101011010010101000: color_data = 12'b111011101110;
20'b00101011010010101001: color_data = 12'b111011101110;
20'b00101011010010101010: color_data = 12'b111011101110;
20'b00101011010011001101: color_data = 12'b111011101110;
20'b00101011010011001110: color_data = 12'b111011101110;
20'b00101011010011001111: color_data = 12'b111011101110;
20'b00101011010011010000: color_data = 12'b111011101110;
20'b00101011010011010001: color_data = 12'b111011101110;
20'b00101011010011010010: color_data = 12'b111011101110;
20'b00101011010011010011: color_data = 12'b111011101110;
20'b00101011010011010100: color_data = 12'b111011101110;
20'b00101011010011010101: color_data = 12'b111011101110;
20'b00101011010011010110: color_data = 12'b111011101110;
20'b00101011010011011000: color_data = 12'b111011101110;
20'b00101011010011011001: color_data = 12'b111011101110;
20'b00101011010011011010: color_data = 12'b111011101110;
20'b00101011010011011011: color_data = 12'b111011101110;
20'b00101011010011011100: color_data = 12'b111011101110;
20'b00101011010011011101: color_data = 12'b111011101110;
20'b00101011010011011110: color_data = 12'b111011101110;
20'b00101011010011011111: color_data = 12'b111011101110;
20'b00101011010011100000: color_data = 12'b111011101110;
20'b00101011010011100001: color_data = 12'b111011101110;
20'b00101011010011101110: color_data = 12'b111011101110;
20'b00101011010011101111: color_data = 12'b111011101110;
20'b00101011010011110000: color_data = 12'b111011101110;
20'b00101011010011110001: color_data = 12'b111011101110;
20'b00101011010011110010: color_data = 12'b111011101110;
20'b00101011010011110011: color_data = 12'b111011101110;
20'b00101011010011110100: color_data = 12'b111011101110;
20'b00101011010011110101: color_data = 12'b111011101110;
20'b00101011010011110110: color_data = 12'b111011101110;
20'b00101011010011110111: color_data = 12'b111011101110;
20'b00101011010011111001: color_data = 12'b111011101110;
20'b00101011010011111010: color_data = 12'b111011101110;
20'b00101011010011111011: color_data = 12'b111011101110;
20'b00101011010011111100: color_data = 12'b111011101110;
20'b00101011010011111101: color_data = 12'b111011101110;
20'b00101011010011111110: color_data = 12'b111011101110;
20'b00101011010011111111: color_data = 12'b111011101110;
20'b00101011010100000000: color_data = 12'b111011101110;
20'b00101011010100000001: color_data = 12'b111011101110;
20'b00101011010100000010: color_data = 12'b111011101110;
20'b00101011010100100101: color_data = 12'b111011101110;
20'b00101011010100100110: color_data = 12'b111011101110;
20'b00101011010100100111: color_data = 12'b111011101110;
20'b00101011010100101000: color_data = 12'b111011101110;
20'b00101011010100101001: color_data = 12'b111011101110;
20'b00101011010100101010: color_data = 12'b111011101110;
20'b00101011010100101011: color_data = 12'b111011101110;
20'b00101011010100101100: color_data = 12'b111011101110;
20'b00101011010100101101: color_data = 12'b111011101110;
20'b00101011010100101110: color_data = 12'b111011101110;
20'b00101011010100110000: color_data = 12'b111011101110;
20'b00101011010100110001: color_data = 12'b111011101110;
20'b00101011010100110010: color_data = 12'b111011101110;
20'b00101011010100110011: color_data = 12'b111011101110;
20'b00101011010100110100: color_data = 12'b111011101110;
20'b00101011010100110101: color_data = 12'b111011101110;
20'b00101011010100110110: color_data = 12'b111011101110;
20'b00101011010100110111: color_data = 12'b111011101110;
20'b00101011010100111000: color_data = 12'b111011101110;
20'b00101011010100111001: color_data = 12'b111011101110;
20'b00101011010101000110: color_data = 12'b111011101110;
20'b00101011010101000111: color_data = 12'b111011101110;
20'b00101011010101001000: color_data = 12'b111011101110;
20'b00101011010101001001: color_data = 12'b111011101110;
20'b00101011010101001010: color_data = 12'b111011101110;
20'b00101011010101001011: color_data = 12'b111011101110;
20'b00101011010101001100: color_data = 12'b111011101110;
20'b00101011010101001101: color_data = 12'b111011101110;
20'b00101011010101001110: color_data = 12'b111011101110;
20'b00101011010101001111: color_data = 12'b111011101110;
20'b00101011010101010001: color_data = 12'b111011101110;
20'b00101011010101010010: color_data = 12'b111011101110;
20'b00101011010101010011: color_data = 12'b111011101110;
20'b00101011010101010100: color_data = 12'b111011101110;
20'b00101011010101010101: color_data = 12'b111011101110;
20'b00101011010101010110: color_data = 12'b111011101110;
20'b00101011010101010111: color_data = 12'b111011101110;
20'b00101011010101011000: color_data = 12'b111011101110;
20'b00101011010101011001: color_data = 12'b111011101110;
20'b00101011010101011010: color_data = 12'b111011101110;
20'b00101011010101111101: color_data = 12'b111011101110;
20'b00101011010101111110: color_data = 12'b111011101110;
20'b00101011010101111111: color_data = 12'b111011101110;
20'b00101011010110000000: color_data = 12'b111011101110;
20'b00101011010110000001: color_data = 12'b111011101110;
20'b00101011010110000010: color_data = 12'b111011101110;
20'b00101011010110000011: color_data = 12'b111011101110;
20'b00101011010110000100: color_data = 12'b111011101110;
20'b00101011010110000101: color_data = 12'b111011101110;
20'b00101011010110000110: color_data = 12'b111011101110;
20'b00101011010110001000: color_data = 12'b111011101110;
20'b00101011010110001001: color_data = 12'b111011101110;
20'b00101011010110001010: color_data = 12'b111011101110;
20'b00101011010110001011: color_data = 12'b111011101110;
20'b00101011010110001100: color_data = 12'b111011101110;
20'b00101011010110001101: color_data = 12'b111011101110;
20'b00101011010110001110: color_data = 12'b111011101110;
20'b00101011010110001111: color_data = 12'b111011101110;
20'b00101011010110010000: color_data = 12'b111011101110;
20'b00101011010110010001: color_data = 12'b111011101110;
20'b00101011010110011110: color_data = 12'b111011101110;
20'b00101011010110011111: color_data = 12'b111011101110;
20'b00101011010110100000: color_data = 12'b111011101110;
20'b00101011010110100001: color_data = 12'b111011101110;
20'b00101011010110100010: color_data = 12'b111011101110;
20'b00101011010110100011: color_data = 12'b111011101110;
20'b00101011010110100100: color_data = 12'b111011101110;
20'b00101011010110100101: color_data = 12'b111011101110;
20'b00101011010110100110: color_data = 12'b111011101110;
20'b00101011010110100111: color_data = 12'b111011101110;
20'b00101011010110101001: color_data = 12'b111011101110;
20'b00101011010110101010: color_data = 12'b111011101110;
20'b00101011010110101011: color_data = 12'b111011101110;
20'b00101011010110101100: color_data = 12'b111011101110;
20'b00101011010110101101: color_data = 12'b111011101110;
20'b00101011010110101110: color_data = 12'b111011101110;
20'b00101011010110101111: color_data = 12'b111011101110;
20'b00101011010110110000: color_data = 12'b111011101110;
20'b00101011010110110001: color_data = 12'b111011101110;
20'b00101011010110110010: color_data = 12'b111011101110;
20'b00101011100010010110: color_data = 12'b111011101110;
20'b00101011100010010111: color_data = 12'b111011101110;
20'b00101011100010011000: color_data = 12'b111011101110;
20'b00101011100010011001: color_data = 12'b111011101110;
20'b00101011100010011010: color_data = 12'b111011101110;
20'b00101011100010011011: color_data = 12'b111011101110;
20'b00101011100010011100: color_data = 12'b111011101110;
20'b00101011100010011101: color_data = 12'b111011101110;
20'b00101011100010011110: color_data = 12'b111011101110;
20'b00101011100010011111: color_data = 12'b111011101110;
20'b00101011100010100001: color_data = 12'b111011101110;
20'b00101011100010100010: color_data = 12'b111011101110;
20'b00101011100010100011: color_data = 12'b111011101110;
20'b00101011100010100100: color_data = 12'b111011101110;
20'b00101011100010100101: color_data = 12'b111011101110;
20'b00101011100010100110: color_data = 12'b111011101110;
20'b00101011100010100111: color_data = 12'b111011101110;
20'b00101011100010101000: color_data = 12'b111011101110;
20'b00101011100010101001: color_data = 12'b111011101110;
20'b00101011100010101010: color_data = 12'b111011101110;
20'b00101011100011001101: color_data = 12'b111011101110;
20'b00101011100011001110: color_data = 12'b111011101110;
20'b00101011100011001111: color_data = 12'b111011101110;
20'b00101011100011010000: color_data = 12'b111011101110;
20'b00101011100011010001: color_data = 12'b111011101110;
20'b00101011100011010010: color_data = 12'b111011101110;
20'b00101011100011010011: color_data = 12'b111011101110;
20'b00101011100011010100: color_data = 12'b111011101110;
20'b00101011100011010101: color_data = 12'b111011101110;
20'b00101011100011010110: color_data = 12'b111011101110;
20'b00101011100011011000: color_data = 12'b111011101110;
20'b00101011100011011001: color_data = 12'b111011101110;
20'b00101011100011011010: color_data = 12'b111011101110;
20'b00101011100011011011: color_data = 12'b111011101110;
20'b00101011100011011100: color_data = 12'b111011101110;
20'b00101011100011011101: color_data = 12'b111011101110;
20'b00101011100011011110: color_data = 12'b111011101110;
20'b00101011100011011111: color_data = 12'b111011101110;
20'b00101011100011100000: color_data = 12'b111011101110;
20'b00101011100011100001: color_data = 12'b111011101110;
20'b00101011100011101110: color_data = 12'b111011101110;
20'b00101011100011101111: color_data = 12'b111011101110;
20'b00101011100011110000: color_data = 12'b111011101110;
20'b00101011100011110001: color_data = 12'b111011101110;
20'b00101011100011110010: color_data = 12'b111011101110;
20'b00101011100011110011: color_data = 12'b111011101110;
20'b00101011100011110100: color_data = 12'b111011101110;
20'b00101011100011110101: color_data = 12'b111011101110;
20'b00101011100011110110: color_data = 12'b111011101110;
20'b00101011100011110111: color_data = 12'b111011101110;
20'b00101011100011111001: color_data = 12'b111011101110;
20'b00101011100011111010: color_data = 12'b111011101110;
20'b00101011100011111011: color_data = 12'b111011101110;
20'b00101011100011111100: color_data = 12'b111011101110;
20'b00101011100011111101: color_data = 12'b111011101110;
20'b00101011100011111110: color_data = 12'b111011101110;
20'b00101011100011111111: color_data = 12'b111011101110;
20'b00101011100100000000: color_data = 12'b111011101110;
20'b00101011100100000001: color_data = 12'b111011101110;
20'b00101011100100000010: color_data = 12'b111011101110;
20'b00101011100100100101: color_data = 12'b111011101110;
20'b00101011100100100110: color_data = 12'b111011101110;
20'b00101011100100100111: color_data = 12'b111011101110;
20'b00101011100100101000: color_data = 12'b111011101110;
20'b00101011100100101001: color_data = 12'b111011101110;
20'b00101011100100101010: color_data = 12'b111011101110;
20'b00101011100100101011: color_data = 12'b111011101110;
20'b00101011100100101100: color_data = 12'b111011101110;
20'b00101011100100101101: color_data = 12'b111011101110;
20'b00101011100100101110: color_data = 12'b111011101110;
20'b00101011100100110000: color_data = 12'b111011101110;
20'b00101011100100110001: color_data = 12'b111011101110;
20'b00101011100100110010: color_data = 12'b111011101110;
20'b00101011100100110011: color_data = 12'b111011101110;
20'b00101011100100110100: color_data = 12'b111011101110;
20'b00101011100100110101: color_data = 12'b111011101110;
20'b00101011100100110110: color_data = 12'b111011101110;
20'b00101011100100110111: color_data = 12'b111011101110;
20'b00101011100100111000: color_data = 12'b111011101110;
20'b00101011100100111001: color_data = 12'b111011101110;
20'b00101011100101000110: color_data = 12'b111011101110;
20'b00101011100101000111: color_data = 12'b111011101110;
20'b00101011100101001000: color_data = 12'b111011101110;
20'b00101011100101001001: color_data = 12'b111011101110;
20'b00101011100101001010: color_data = 12'b111011101110;
20'b00101011100101001011: color_data = 12'b111011101110;
20'b00101011100101001100: color_data = 12'b111011101110;
20'b00101011100101001101: color_data = 12'b111011101110;
20'b00101011100101001110: color_data = 12'b111011101110;
20'b00101011100101001111: color_data = 12'b111011101110;
20'b00101011100101010001: color_data = 12'b111011101110;
20'b00101011100101010010: color_data = 12'b111011101110;
20'b00101011100101010011: color_data = 12'b111011101110;
20'b00101011100101010100: color_data = 12'b111011101110;
20'b00101011100101010101: color_data = 12'b111011101110;
20'b00101011100101010110: color_data = 12'b111011101110;
20'b00101011100101010111: color_data = 12'b111011101110;
20'b00101011100101011000: color_data = 12'b111011101110;
20'b00101011100101011001: color_data = 12'b111011101110;
20'b00101011100101011010: color_data = 12'b111011101110;
20'b00101011100101111101: color_data = 12'b111011101110;
20'b00101011100101111110: color_data = 12'b111011101110;
20'b00101011100101111111: color_data = 12'b111011101110;
20'b00101011100110000000: color_data = 12'b111011101110;
20'b00101011100110000001: color_data = 12'b111011101110;
20'b00101011100110000010: color_data = 12'b111011101110;
20'b00101011100110000011: color_data = 12'b111011101110;
20'b00101011100110000100: color_data = 12'b111011101110;
20'b00101011100110000101: color_data = 12'b111011101110;
20'b00101011100110000110: color_data = 12'b111011101110;
20'b00101011100110001000: color_data = 12'b111011101110;
20'b00101011100110001001: color_data = 12'b111011101110;
20'b00101011100110001010: color_data = 12'b111011101110;
20'b00101011100110001011: color_data = 12'b111011101110;
20'b00101011100110001100: color_data = 12'b111011101110;
20'b00101011100110001101: color_data = 12'b111011101110;
20'b00101011100110001110: color_data = 12'b111011101110;
20'b00101011100110001111: color_data = 12'b111011101110;
20'b00101011100110010000: color_data = 12'b111011101110;
20'b00101011100110010001: color_data = 12'b111011101110;
20'b00101011100110011110: color_data = 12'b111011101110;
20'b00101011100110011111: color_data = 12'b111011101110;
20'b00101011100110100000: color_data = 12'b111011101110;
20'b00101011100110100001: color_data = 12'b111011101110;
20'b00101011100110100010: color_data = 12'b111011101110;
20'b00101011100110100011: color_data = 12'b111011101110;
20'b00101011100110100100: color_data = 12'b111011101110;
20'b00101011100110100101: color_data = 12'b111011101110;
20'b00101011100110100110: color_data = 12'b111011101110;
20'b00101011100110100111: color_data = 12'b111011101110;
20'b00101011100110101001: color_data = 12'b111011101110;
20'b00101011100110101010: color_data = 12'b111011101110;
20'b00101011100110101011: color_data = 12'b111011101110;
20'b00101011100110101100: color_data = 12'b111011101110;
20'b00101011100110101101: color_data = 12'b111011101110;
20'b00101011100110101110: color_data = 12'b111011101110;
20'b00101011100110101111: color_data = 12'b111011101110;
20'b00101011100110110000: color_data = 12'b111011101110;
20'b00101011100110110001: color_data = 12'b111011101110;
20'b00101011100110110010: color_data = 12'b111011101110;
20'b00101011110010010110: color_data = 12'b111011101110;
20'b00101011110010010111: color_data = 12'b111011101110;
20'b00101011110010011000: color_data = 12'b111011101110;
20'b00101011110010011001: color_data = 12'b111011101110;
20'b00101011110010011010: color_data = 12'b111011101110;
20'b00101011110010011011: color_data = 12'b111011101110;
20'b00101011110010011100: color_data = 12'b111011101110;
20'b00101011110010011101: color_data = 12'b111011101110;
20'b00101011110010011110: color_data = 12'b111011101110;
20'b00101011110010011111: color_data = 12'b111011101110;
20'b00101011110010100001: color_data = 12'b111011101110;
20'b00101011110010100010: color_data = 12'b111011101110;
20'b00101011110010100011: color_data = 12'b111011101110;
20'b00101011110010100100: color_data = 12'b111011101110;
20'b00101011110010100101: color_data = 12'b111011101110;
20'b00101011110010100110: color_data = 12'b111011101110;
20'b00101011110010100111: color_data = 12'b111011101110;
20'b00101011110010101000: color_data = 12'b111011101110;
20'b00101011110010101001: color_data = 12'b111011101110;
20'b00101011110010101010: color_data = 12'b111011101110;
20'b00101011110011001101: color_data = 12'b111011101110;
20'b00101011110011001110: color_data = 12'b111011101110;
20'b00101011110011001111: color_data = 12'b111011101110;
20'b00101011110011010000: color_data = 12'b111011101110;
20'b00101011110011010001: color_data = 12'b111011101110;
20'b00101011110011010010: color_data = 12'b111011101110;
20'b00101011110011010011: color_data = 12'b111011101110;
20'b00101011110011010100: color_data = 12'b111011101110;
20'b00101011110011010101: color_data = 12'b111011101110;
20'b00101011110011010110: color_data = 12'b111011101110;
20'b00101011110011011000: color_data = 12'b111011101110;
20'b00101011110011011001: color_data = 12'b111011101110;
20'b00101011110011011010: color_data = 12'b111011101110;
20'b00101011110011011011: color_data = 12'b111011101110;
20'b00101011110011011100: color_data = 12'b111011101110;
20'b00101011110011011101: color_data = 12'b111011101110;
20'b00101011110011011110: color_data = 12'b111011101110;
20'b00101011110011011111: color_data = 12'b111011101110;
20'b00101011110011100000: color_data = 12'b111011101110;
20'b00101011110011100001: color_data = 12'b111011101110;
20'b00101011110011101110: color_data = 12'b111011101110;
20'b00101011110011101111: color_data = 12'b111011101110;
20'b00101011110011110000: color_data = 12'b111011101110;
20'b00101011110011110001: color_data = 12'b111011101110;
20'b00101011110011110010: color_data = 12'b111011101110;
20'b00101011110011110011: color_data = 12'b111011101110;
20'b00101011110011110100: color_data = 12'b111011101110;
20'b00101011110011110101: color_data = 12'b111011101110;
20'b00101011110011110110: color_data = 12'b111011101110;
20'b00101011110011110111: color_data = 12'b111011101110;
20'b00101011110011111001: color_data = 12'b111011101110;
20'b00101011110011111010: color_data = 12'b111011101110;
20'b00101011110011111011: color_data = 12'b111011101110;
20'b00101011110011111100: color_data = 12'b111011101110;
20'b00101011110011111101: color_data = 12'b111011101110;
20'b00101011110011111110: color_data = 12'b111011101110;
20'b00101011110011111111: color_data = 12'b111011101110;
20'b00101011110100000000: color_data = 12'b111011101110;
20'b00101011110100000001: color_data = 12'b111011101110;
20'b00101011110100000010: color_data = 12'b111011101110;
20'b00101011110100100101: color_data = 12'b111011101110;
20'b00101011110100100110: color_data = 12'b111011101110;
20'b00101011110100100111: color_data = 12'b111011101110;
20'b00101011110100101000: color_data = 12'b111011101110;
20'b00101011110100101001: color_data = 12'b111011101110;
20'b00101011110100101010: color_data = 12'b111011101110;
20'b00101011110100101011: color_data = 12'b111011101110;
20'b00101011110100101100: color_data = 12'b111011101110;
20'b00101011110100101101: color_data = 12'b111011101110;
20'b00101011110100101110: color_data = 12'b111011101110;
20'b00101011110100110000: color_data = 12'b111011101110;
20'b00101011110100110001: color_data = 12'b111011101110;
20'b00101011110100110010: color_data = 12'b111011101110;
20'b00101011110100110011: color_data = 12'b111011101110;
20'b00101011110100110100: color_data = 12'b111011101110;
20'b00101011110100110101: color_data = 12'b111011101110;
20'b00101011110100110110: color_data = 12'b111011101110;
20'b00101011110100110111: color_data = 12'b111011101110;
20'b00101011110100111000: color_data = 12'b111011101110;
20'b00101011110100111001: color_data = 12'b111011101110;
20'b00101011110101000110: color_data = 12'b111011101110;
20'b00101011110101000111: color_data = 12'b111011101110;
20'b00101011110101001000: color_data = 12'b111011101110;
20'b00101011110101001001: color_data = 12'b111011101110;
20'b00101011110101001010: color_data = 12'b111011101110;
20'b00101011110101001011: color_data = 12'b111011101110;
20'b00101011110101001100: color_data = 12'b111011101110;
20'b00101011110101001101: color_data = 12'b111011101110;
20'b00101011110101001110: color_data = 12'b111011101110;
20'b00101011110101001111: color_data = 12'b111011101110;
20'b00101011110101010001: color_data = 12'b111011101110;
20'b00101011110101010010: color_data = 12'b111011101110;
20'b00101011110101010011: color_data = 12'b111011101110;
20'b00101011110101010100: color_data = 12'b111011101110;
20'b00101011110101010101: color_data = 12'b111011101110;
20'b00101011110101010110: color_data = 12'b111011101110;
20'b00101011110101010111: color_data = 12'b111011101110;
20'b00101011110101011000: color_data = 12'b111011101110;
20'b00101011110101011001: color_data = 12'b111011101110;
20'b00101011110101011010: color_data = 12'b111011101110;
20'b00101011110101111101: color_data = 12'b111011101110;
20'b00101011110101111110: color_data = 12'b111011101110;
20'b00101011110101111111: color_data = 12'b111011101110;
20'b00101011110110000000: color_data = 12'b111011101110;
20'b00101011110110000001: color_data = 12'b111011101110;
20'b00101011110110000010: color_data = 12'b111011101110;
20'b00101011110110000011: color_data = 12'b111011101110;
20'b00101011110110000100: color_data = 12'b111011101110;
20'b00101011110110000101: color_data = 12'b111011101110;
20'b00101011110110000110: color_data = 12'b111011101110;
20'b00101011110110001000: color_data = 12'b111011101110;
20'b00101011110110001001: color_data = 12'b111011101110;
20'b00101011110110001010: color_data = 12'b111011101110;
20'b00101011110110001011: color_data = 12'b111011101110;
20'b00101011110110001100: color_data = 12'b111011101110;
20'b00101011110110001101: color_data = 12'b111011101110;
20'b00101011110110001110: color_data = 12'b111011101110;
20'b00101011110110001111: color_data = 12'b111011101110;
20'b00101011110110010000: color_data = 12'b111011101110;
20'b00101011110110010001: color_data = 12'b111011101110;
20'b00101011110110011110: color_data = 12'b111011101110;
20'b00101011110110011111: color_data = 12'b111011101110;
20'b00101011110110100000: color_data = 12'b111011101110;
20'b00101011110110100001: color_data = 12'b111011101110;
20'b00101011110110100010: color_data = 12'b111011101110;
20'b00101011110110100011: color_data = 12'b111011101110;
20'b00101011110110100100: color_data = 12'b111011101110;
20'b00101011110110100101: color_data = 12'b111011101110;
20'b00101011110110100110: color_data = 12'b111011101110;
20'b00101011110110100111: color_data = 12'b111011101110;
20'b00101011110110101001: color_data = 12'b111011101110;
20'b00101011110110101010: color_data = 12'b111011101110;
20'b00101011110110101011: color_data = 12'b111011101110;
20'b00101011110110101100: color_data = 12'b111011101110;
20'b00101011110110101101: color_data = 12'b111011101110;
20'b00101011110110101110: color_data = 12'b111011101110;
20'b00101011110110101111: color_data = 12'b111011101110;
20'b00101011110110110000: color_data = 12'b111011101110;
20'b00101011110110110001: color_data = 12'b111011101110;
20'b00101011110110110010: color_data = 12'b111011101110;
20'b00101100010010010110: color_data = 12'b111011101110;
20'b00101100010010010111: color_data = 12'b111011101110;
20'b00101100010010011000: color_data = 12'b111011101110;
20'b00101100010010011001: color_data = 12'b111011101110;
20'b00101100010010011010: color_data = 12'b111011101110;
20'b00101100010010011011: color_data = 12'b111011101110;
20'b00101100010010011100: color_data = 12'b111011101110;
20'b00101100010010011101: color_data = 12'b111011101110;
20'b00101100010010011110: color_data = 12'b111011101110;
20'b00101100010010011111: color_data = 12'b111011101110;
20'b00101100010010100001: color_data = 12'b111011101110;
20'b00101100010010100010: color_data = 12'b111011101110;
20'b00101100010010100011: color_data = 12'b111011101110;
20'b00101100010010100100: color_data = 12'b111011101110;
20'b00101100010010100101: color_data = 12'b111011101110;
20'b00101100010010100110: color_data = 12'b111011101110;
20'b00101100010010100111: color_data = 12'b111011101110;
20'b00101100010010101000: color_data = 12'b111011101110;
20'b00101100010010101001: color_data = 12'b111011101110;
20'b00101100010010101010: color_data = 12'b111011101110;
20'b00101100010010101100: color_data = 12'b111011101110;
20'b00101100010010101101: color_data = 12'b111011101110;
20'b00101100010010101110: color_data = 12'b111011101110;
20'b00101100010010101111: color_data = 12'b111011101110;
20'b00101100010010110000: color_data = 12'b111011101110;
20'b00101100010010110001: color_data = 12'b111011101110;
20'b00101100010010110010: color_data = 12'b111011101110;
20'b00101100010010110011: color_data = 12'b111011101110;
20'b00101100010010110100: color_data = 12'b111011101110;
20'b00101100010010110101: color_data = 12'b111011101110;
20'b00101100010010110111: color_data = 12'b111011101110;
20'b00101100010010111000: color_data = 12'b111011101110;
20'b00101100010010111001: color_data = 12'b111011101110;
20'b00101100010010111010: color_data = 12'b111011101110;
20'b00101100010010111011: color_data = 12'b111011101110;
20'b00101100010010111100: color_data = 12'b111011101110;
20'b00101100010010111101: color_data = 12'b111011101110;
20'b00101100010010111110: color_data = 12'b111011101110;
20'b00101100010010111111: color_data = 12'b111011101110;
20'b00101100010011000000: color_data = 12'b111011101110;
20'b00101100010011000010: color_data = 12'b111011101110;
20'b00101100010011000011: color_data = 12'b111011101110;
20'b00101100010011000100: color_data = 12'b111011101110;
20'b00101100010011000101: color_data = 12'b111011101110;
20'b00101100010011000110: color_data = 12'b111011101110;
20'b00101100010011000111: color_data = 12'b111011101110;
20'b00101100010011001000: color_data = 12'b111011101110;
20'b00101100010011001001: color_data = 12'b111011101110;
20'b00101100010011001010: color_data = 12'b111011101110;
20'b00101100010011001011: color_data = 12'b111011101110;
20'b00101100010011001101: color_data = 12'b111011101110;
20'b00101100010011001110: color_data = 12'b111011101110;
20'b00101100010011001111: color_data = 12'b111011101110;
20'b00101100010011010000: color_data = 12'b111011101110;
20'b00101100010011010001: color_data = 12'b111011101110;
20'b00101100010011010010: color_data = 12'b111011101110;
20'b00101100010011010011: color_data = 12'b111011101110;
20'b00101100010011010100: color_data = 12'b111011101110;
20'b00101100010011010101: color_data = 12'b111011101110;
20'b00101100010011010110: color_data = 12'b111011101110;
20'b00101100010011011000: color_data = 12'b111011101110;
20'b00101100010011011001: color_data = 12'b111011101110;
20'b00101100010011011010: color_data = 12'b111011101110;
20'b00101100010011011011: color_data = 12'b111011101110;
20'b00101100010011011100: color_data = 12'b111011101110;
20'b00101100010011011101: color_data = 12'b111011101110;
20'b00101100010011011110: color_data = 12'b111011101110;
20'b00101100010011011111: color_data = 12'b111011101110;
20'b00101100010011100000: color_data = 12'b111011101110;
20'b00101100010011100001: color_data = 12'b111011101110;
20'b00101100010011101110: color_data = 12'b111011101110;
20'b00101100010011101111: color_data = 12'b111011101110;
20'b00101100010011110000: color_data = 12'b111011101110;
20'b00101100010011110001: color_data = 12'b111011101110;
20'b00101100010011110010: color_data = 12'b111011101110;
20'b00101100010011110011: color_data = 12'b111011101110;
20'b00101100010011110100: color_data = 12'b111011101110;
20'b00101100010011110101: color_data = 12'b111011101110;
20'b00101100010011110110: color_data = 12'b111011101110;
20'b00101100010011110111: color_data = 12'b111011101110;
20'b00101100010011111001: color_data = 12'b111011101110;
20'b00101100010011111010: color_data = 12'b111011101110;
20'b00101100010011111011: color_data = 12'b111011101110;
20'b00101100010011111100: color_data = 12'b111011101110;
20'b00101100010011111101: color_data = 12'b111011101110;
20'b00101100010011111110: color_data = 12'b111011101110;
20'b00101100010011111111: color_data = 12'b111011101110;
20'b00101100010100000000: color_data = 12'b111011101110;
20'b00101100010100000001: color_data = 12'b111011101110;
20'b00101100010100000010: color_data = 12'b111011101110;
20'b00101100010100100101: color_data = 12'b111011101110;
20'b00101100010100100110: color_data = 12'b111011101110;
20'b00101100010100100111: color_data = 12'b111011101110;
20'b00101100010100101000: color_data = 12'b111011101110;
20'b00101100010100101001: color_data = 12'b111011101110;
20'b00101100010100101010: color_data = 12'b111011101110;
20'b00101100010100101011: color_data = 12'b111011101110;
20'b00101100010100101100: color_data = 12'b111011101110;
20'b00101100010100101101: color_data = 12'b111011101110;
20'b00101100010100101110: color_data = 12'b111011101110;
20'b00101100010100110000: color_data = 12'b111011101110;
20'b00101100010100110001: color_data = 12'b111011101110;
20'b00101100010100110010: color_data = 12'b111011101110;
20'b00101100010100110011: color_data = 12'b111011101110;
20'b00101100010100110100: color_data = 12'b111011101110;
20'b00101100010100110101: color_data = 12'b111011101110;
20'b00101100010100110110: color_data = 12'b111011101110;
20'b00101100010100110111: color_data = 12'b111011101110;
20'b00101100010100111000: color_data = 12'b111011101110;
20'b00101100010100111001: color_data = 12'b111011101110;
20'b00101100010101000110: color_data = 12'b111011101110;
20'b00101100010101000111: color_data = 12'b111011101110;
20'b00101100010101001000: color_data = 12'b111011101110;
20'b00101100010101001001: color_data = 12'b111011101110;
20'b00101100010101001010: color_data = 12'b111011101110;
20'b00101100010101001011: color_data = 12'b111011101110;
20'b00101100010101001100: color_data = 12'b111011101110;
20'b00101100010101001101: color_data = 12'b111011101110;
20'b00101100010101001110: color_data = 12'b111011101110;
20'b00101100010101001111: color_data = 12'b111011101110;
20'b00101100010101010001: color_data = 12'b111011101110;
20'b00101100010101010010: color_data = 12'b111011101110;
20'b00101100010101010011: color_data = 12'b111011101110;
20'b00101100010101010100: color_data = 12'b111011101110;
20'b00101100010101010101: color_data = 12'b111011101110;
20'b00101100010101010110: color_data = 12'b111011101110;
20'b00101100010101010111: color_data = 12'b111011101110;
20'b00101100010101011000: color_data = 12'b111011101110;
20'b00101100010101011001: color_data = 12'b111011101110;
20'b00101100010101011010: color_data = 12'b111011101110;
20'b00101100010101111101: color_data = 12'b111011101110;
20'b00101100010101111110: color_data = 12'b111011101110;
20'b00101100010101111111: color_data = 12'b111011101110;
20'b00101100010110000000: color_data = 12'b111011101110;
20'b00101100010110000001: color_data = 12'b111011101110;
20'b00101100010110000010: color_data = 12'b111011101110;
20'b00101100010110000011: color_data = 12'b111011101110;
20'b00101100010110000100: color_data = 12'b111011101110;
20'b00101100010110000101: color_data = 12'b111011101110;
20'b00101100010110000110: color_data = 12'b111011101110;
20'b00101100010110001000: color_data = 12'b111011101110;
20'b00101100010110001001: color_data = 12'b111011101110;
20'b00101100010110001010: color_data = 12'b111011101110;
20'b00101100010110001011: color_data = 12'b111011101110;
20'b00101100010110001100: color_data = 12'b111011101110;
20'b00101100010110001101: color_data = 12'b111011101110;
20'b00101100010110001110: color_data = 12'b111011101110;
20'b00101100010110001111: color_data = 12'b111011101110;
20'b00101100010110010000: color_data = 12'b111011101110;
20'b00101100010110010001: color_data = 12'b111011101110;
20'b00101100010110011110: color_data = 12'b111011101110;
20'b00101100010110011111: color_data = 12'b111011101110;
20'b00101100010110100000: color_data = 12'b111011101110;
20'b00101100010110100001: color_data = 12'b111011101110;
20'b00101100010110100010: color_data = 12'b111011101110;
20'b00101100010110100011: color_data = 12'b111011101110;
20'b00101100010110100100: color_data = 12'b111011101110;
20'b00101100010110100101: color_data = 12'b111011101110;
20'b00101100010110100110: color_data = 12'b111011101110;
20'b00101100010110100111: color_data = 12'b111011101110;
20'b00101100010110101001: color_data = 12'b111011101110;
20'b00101100010110101010: color_data = 12'b111011101110;
20'b00101100010110101011: color_data = 12'b111011101110;
20'b00101100010110101100: color_data = 12'b111011101110;
20'b00101100010110101101: color_data = 12'b111011101110;
20'b00101100010110101110: color_data = 12'b111011101110;
20'b00101100010110101111: color_data = 12'b111011101110;
20'b00101100010110110000: color_data = 12'b111011101110;
20'b00101100010110110001: color_data = 12'b111011101110;
20'b00101100010110110010: color_data = 12'b111011101110;
20'b00101100010110110100: color_data = 12'b111011101110;
20'b00101100010110110101: color_data = 12'b111011101110;
20'b00101100010110110110: color_data = 12'b111011101110;
20'b00101100010110110111: color_data = 12'b111011101110;
20'b00101100010110111000: color_data = 12'b111011101110;
20'b00101100010110111001: color_data = 12'b111011101110;
20'b00101100010110111010: color_data = 12'b111011101110;
20'b00101100010110111011: color_data = 12'b111011101110;
20'b00101100010110111100: color_data = 12'b111011101110;
20'b00101100010110111101: color_data = 12'b111011101110;
20'b00101100010110111111: color_data = 12'b111011101110;
20'b00101100010111000000: color_data = 12'b111011101110;
20'b00101100010111000001: color_data = 12'b111011101110;
20'b00101100010111000010: color_data = 12'b111011101110;
20'b00101100010111000011: color_data = 12'b111011101110;
20'b00101100010111000100: color_data = 12'b111011101110;
20'b00101100010111000101: color_data = 12'b111011101110;
20'b00101100010111000110: color_data = 12'b111011101110;
20'b00101100010111000111: color_data = 12'b111011101110;
20'b00101100010111001000: color_data = 12'b111011101110;
20'b00101100010111001010: color_data = 12'b111011101110;
20'b00101100010111001011: color_data = 12'b111011101110;
20'b00101100010111001100: color_data = 12'b111011101110;
20'b00101100010111001101: color_data = 12'b111011101110;
20'b00101100010111001110: color_data = 12'b111011101110;
20'b00101100010111001111: color_data = 12'b111011101110;
20'b00101100010111010000: color_data = 12'b111011101110;
20'b00101100010111010001: color_data = 12'b111011101110;
20'b00101100010111010010: color_data = 12'b111011101110;
20'b00101100010111010011: color_data = 12'b111011101110;
20'b00101100010111010101: color_data = 12'b111011101110;
20'b00101100010111010110: color_data = 12'b111011101110;
20'b00101100010111010111: color_data = 12'b111011101110;
20'b00101100010111011000: color_data = 12'b111011101110;
20'b00101100010111011001: color_data = 12'b111011101110;
20'b00101100010111011010: color_data = 12'b111011101110;
20'b00101100010111011011: color_data = 12'b111011101110;
20'b00101100010111011100: color_data = 12'b111011101110;
20'b00101100010111011101: color_data = 12'b111011101110;
20'b00101100010111011110: color_data = 12'b111011101110;
20'b00101100010111100000: color_data = 12'b111011101110;
20'b00101100010111100001: color_data = 12'b111011101110;
20'b00101100010111100010: color_data = 12'b111011101110;
20'b00101100010111100011: color_data = 12'b111011101110;
20'b00101100010111100100: color_data = 12'b111011101110;
20'b00101100010111100101: color_data = 12'b111011101110;
20'b00101100010111100110: color_data = 12'b111011101110;
20'b00101100010111100111: color_data = 12'b111011101110;
20'b00101100010111101000: color_data = 12'b111011101110;
20'b00101100010111101001: color_data = 12'b111011101110;
20'b00101100100010010110: color_data = 12'b111011101110;
20'b00101100100010010111: color_data = 12'b111011101110;
20'b00101100100010011000: color_data = 12'b111011101110;
20'b00101100100010011001: color_data = 12'b111011101110;
20'b00101100100010011010: color_data = 12'b111011101110;
20'b00101100100010011011: color_data = 12'b111011101110;
20'b00101100100010011100: color_data = 12'b111011101110;
20'b00101100100010011101: color_data = 12'b111011101110;
20'b00101100100010011110: color_data = 12'b111011101110;
20'b00101100100010011111: color_data = 12'b111011101110;
20'b00101100100010100001: color_data = 12'b111011101110;
20'b00101100100010100010: color_data = 12'b111011101110;
20'b00101100100010100011: color_data = 12'b111011101110;
20'b00101100100010100100: color_data = 12'b111011101110;
20'b00101100100010100101: color_data = 12'b111011101110;
20'b00101100100010100110: color_data = 12'b111011101110;
20'b00101100100010100111: color_data = 12'b111011101110;
20'b00101100100010101000: color_data = 12'b111011101110;
20'b00101100100010101001: color_data = 12'b111011101110;
20'b00101100100010101010: color_data = 12'b111011101110;
20'b00101100100010101100: color_data = 12'b111011101110;
20'b00101100100010101101: color_data = 12'b111011101110;
20'b00101100100010101110: color_data = 12'b111011101110;
20'b00101100100010101111: color_data = 12'b111011101110;
20'b00101100100010110000: color_data = 12'b111011101110;
20'b00101100100010110001: color_data = 12'b111011101110;
20'b00101100100010110010: color_data = 12'b111011101110;
20'b00101100100010110011: color_data = 12'b111011101110;
20'b00101100100010110100: color_data = 12'b111011101110;
20'b00101100100010110101: color_data = 12'b111011101110;
20'b00101100100010110111: color_data = 12'b111011101110;
20'b00101100100010111000: color_data = 12'b111011101110;
20'b00101100100010111001: color_data = 12'b111011101110;
20'b00101100100010111010: color_data = 12'b111011101110;
20'b00101100100010111011: color_data = 12'b111011101110;
20'b00101100100010111100: color_data = 12'b111011101110;
20'b00101100100010111101: color_data = 12'b111011101110;
20'b00101100100010111110: color_data = 12'b111011101110;
20'b00101100100010111111: color_data = 12'b111011101110;
20'b00101100100011000000: color_data = 12'b111011101110;
20'b00101100100011000010: color_data = 12'b111011101110;
20'b00101100100011000011: color_data = 12'b111011101110;
20'b00101100100011000100: color_data = 12'b111011101110;
20'b00101100100011000101: color_data = 12'b111011101110;
20'b00101100100011000110: color_data = 12'b111011101110;
20'b00101100100011000111: color_data = 12'b111011101110;
20'b00101100100011001000: color_data = 12'b111011101110;
20'b00101100100011001001: color_data = 12'b111011101110;
20'b00101100100011001010: color_data = 12'b111011101110;
20'b00101100100011001011: color_data = 12'b111011101110;
20'b00101100100011001101: color_data = 12'b111011101110;
20'b00101100100011001110: color_data = 12'b111011101110;
20'b00101100100011001111: color_data = 12'b111011101110;
20'b00101100100011010000: color_data = 12'b111011101110;
20'b00101100100011010001: color_data = 12'b111011101110;
20'b00101100100011010010: color_data = 12'b111011101110;
20'b00101100100011010011: color_data = 12'b111011101110;
20'b00101100100011010100: color_data = 12'b111011101110;
20'b00101100100011010101: color_data = 12'b111011101110;
20'b00101100100011010110: color_data = 12'b111011101110;
20'b00101100100011011000: color_data = 12'b111011101110;
20'b00101100100011011001: color_data = 12'b111011101110;
20'b00101100100011011010: color_data = 12'b111011101110;
20'b00101100100011011011: color_data = 12'b111011101110;
20'b00101100100011011100: color_data = 12'b111011101110;
20'b00101100100011011101: color_data = 12'b111011101110;
20'b00101100100011011110: color_data = 12'b111011101110;
20'b00101100100011011111: color_data = 12'b111011101110;
20'b00101100100011100000: color_data = 12'b111011101110;
20'b00101100100011100001: color_data = 12'b111011101110;
20'b00101100100011101110: color_data = 12'b111011101110;
20'b00101100100011101111: color_data = 12'b111011101110;
20'b00101100100011110000: color_data = 12'b111011101110;
20'b00101100100011110001: color_data = 12'b111011101110;
20'b00101100100011110010: color_data = 12'b111011101110;
20'b00101100100011110011: color_data = 12'b111011101110;
20'b00101100100011110100: color_data = 12'b111011101110;
20'b00101100100011110101: color_data = 12'b111011101110;
20'b00101100100011110110: color_data = 12'b111011101110;
20'b00101100100011110111: color_data = 12'b111011101110;
20'b00101100100011111001: color_data = 12'b111011101110;
20'b00101100100011111010: color_data = 12'b111011101110;
20'b00101100100011111011: color_data = 12'b111011101110;
20'b00101100100011111100: color_data = 12'b111011101110;
20'b00101100100011111101: color_data = 12'b111011101110;
20'b00101100100011111110: color_data = 12'b111011101110;
20'b00101100100011111111: color_data = 12'b111011101110;
20'b00101100100100000000: color_data = 12'b111011101110;
20'b00101100100100000001: color_data = 12'b111011101110;
20'b00101100100100000010: color_data = 12'b111011101110;
20'b00101100100100100101: color_data = 12'b111011101110;
20'b00101100100100100110: color_data = 12'b111011101110;
20'b00101100100100100111: color_data = 12'b111011101110;
20'b00101100100100101000: color_data = 12'b111011101110;
20'b00101100100100101001: color_data = 12'b111011101110;
20'b00101100100100101010: color_data = 12'b111011101110;
20'b00101100100100101011: color_data = 12'b111011101110;
20'b00101100100100101100: color_data = 12'b111011101110;
20'b00101100100100101101: color_data = 12'b111011101110;
20'b00101100100100101110: color_data = 12'b111011101110;
20'b00101100100100110000: color_data = 12'b111011101110;
20'b00101100100100110001: color_data = 12'b111011101110;
20'b00101100100100110010: color_data = 12'b111011101110;
20'b00101100100100110011: color_data = 12'b111011101110;
20'b00101100100100110100: color_data = 12'b111011101110;
20'b00101100100100110101: color_data = 12'b111011101110;
20'b00101100100100110110: color_data = 12'b111011101110;
20'b00101100100100110111: color_data = 12'b111011101110;
20'b00101100100100111000: color_data = 12'b111011101110;
20'b00101100100100111001: color_data = 12'b111011101110;
20'b00101100100101000110: color_data = 12'b111011101110;
20'b00101100100101000111: color_data = 12'b111011101110;
20'b00101100100101001000: color_data = 12'b111011101110;
20'b00101100100101001001: color_data = 12'b111011101110;
20'b00101100100101001010: color_data = 12'b111011101110;
20'b00101100100101001011: color_data = 12'b111011101110;
20'b00101100100101001100: color_data = 12'b111011101110;
20'b00101100100101001101: color_data = 12'b111011101110;
20'b00101100100101001110: color_data = 12'b111011101110;
20'b00101100100101001111: color_data = 12'b111011101110;
20'b00101100100101010001: color_data = 12'b111011101110;
20'b00101100100101010010: color_data = 12'b111011101110;
20'b00101100100101010011: color_data = 12'b111011101110;
20'b00101100100101010100: color_data = 12'b111011101110;
20'b00101100100101010101: color_data = 12'b111011101110;
20'b00101100100101010110: color_data = 12'b111011101110;
20'b00101100100101010111: color_data = 12'b111011101110;
20'b00101100100101011000: color_data = 12'b111011101110;
20'b00101100100101011001: color_data = 12'b111011101110;
20'b00101100100101011010: color_data = 12'b111011101110;
20'b00101100100101111101: color_data = 12'b111011101110;
20'b00101100100101111110: color_data = 12'b111011101110;
20'b00101100100101111111: color_data = 12'b111011101110;
20'b00101100100110000000: color_data = 12'b111011101110;
20'b00101100100110000001: color_data = 12'b111011101110;
20'b00101100100110000010: color_data = 12'b111011101110;
20'b00101100100110000011: color_data = 12'b111011101110;
20'b00101100100110000100: color_data = 12'b111011101110;
20'b00101100100110000101: color_data = 12'b111011101110;
20'b00101100100110000110: color_data = 12'b111011101110;
20'b00101100100110001000: color_data = 12'b111011101110;
20'b00101100100110001001: color_data = 12'b111011101110;
20'b00101100100110001010: color_data = 12'b111011101110;
20'b00101100100110001011: color_data = 12'b111011101110;
20'b00101100100110001100: color_data = 12'b111011101110;
20'b00101100100110001101: color_data = 12'b111011101110;
20'b00101100100110001110: color_data = 12'b111011101110;
20'b00101100100110001111: color_data = 12'b111011101110;
20'b00101100100110010000: color_data = 12'b111011101110;
20'b00101100100110010001: color_data = 12'b111011101110;
20'b00101100100110011110: color_data = 12'b111011101110;
20'b00101100100110011111: color_data = 12'b111011101110;
20'b00101100100110100000: color_data = 12'b111011101110;
20'b00101100100110100001: color_data = 12'b111011101110;
20'b00101100100110100010: color_data = 12'b111011101110;
20'b00101100100110100011: color_data = 12'b111011101110;
20'b00101100100110100100: color_data = 12'b111011101110;
20'b00101100100110100101: color_data = 12'b111011101110;
20'b00101100100110100110: color_data = 12'b111011101110;
20'b00101100100110100111: color_data = 12'b111011101110;
20'b00101100100110101001: color_data = 12'b111011101110;
20'b00101100100110101010: color_data = 12'b111011101110;
20'b00101100100110101011: color_data = 12'b111011101110;
20'b00101100100110101100: color_data = 12'b111011101110;
20'b00101100100110101101: color_data = 12'b111011101110;
20'b00101100100110101110: color_data = 12'b111011101110;
20'b00101100100110101111: color_data = 12'b111011101110;
20'b00101100100110110000: color_data = 12'b111011101110;
20'b00101100100110110001: color_data = 12'b111011101110;
20'b00101100100110110010: color_data = 12'b111011101110;
20'b00101100100110110100: color_data = 12'b111011101110;
20'b00101100100110110101: color_data = 12'b111011101110;
20'b00101100100110110110: color_data = 12'b111011101110;
20'b00101100100110110111: color_data = 12'b111011101110;
20'b00101100100110111000: color_data = 12'b111011101110;
20'b00101100100110111001: color_data = 12'b111011101110;
20'b00101100100110111010: color_data = 12'b111011101110;
20'b00101100100110111011: color_data = 12'b111011101110;
20'b00101100100110111100: color_data = 12'b111011101110;
20'b00101100100110111101: color_data = 12'b111011101110;
20'b00101100100110111111: color_data = 12'b111011101110;
20'b00101100100111000000: color_data = 12'b111011101110;
20'b00101100100111000001: color_data = 12'b111011101110;
20'b00101100100111000010: color_data = 12'b111011101110;
20'b00101100100111000011: color_data = 12'b111011101110;
20'b00101100100111000100: color_data = 12'b111011101110;
20'b00101100100111000101: color_data = 12'b111011101110;
20'b00101100100111000110: color_data = 12'b111011101110;
20'b00101100100111000111: color_data = 12'b111011101110;
20'b00101100100111001000: color_data = 12'b111011101110;
20'b00101100100111001010: color_data = 12'b111011101110;
20'b00101100100111001011: color_data = 12'b111011101110;
20'b00101100100111001100: color_data = 12'b111011101110;
20'b00101100100111001101: color_data = 12'b111011101110;
20'b00101100100111001110: color_data = 12'b111011101110;
20'b00101100100111001111: color_data = 12'b111011101110;
20'b00101100100111010000: color_data = 12'b111011101110;
20'b00101100100111010001: color_data = 12'b111011101110;
20'b00101100100111010010: color_data = 12'b111011101110;
20'b00101100100111010011: color_data = 12'b111011101110;
20'b00101100100111010101: color_data = 12'b111011101110;
20'b00101100100111010110: color_data = 12'b111011101110;
20'b00101100100111010111: color_data = 12'b111011101110;
20'b00101100100111011000: color_data = 12'b111011101110;
20'b00101100100111011001: color_data = 12'b111011101110;
20'b00101100100111011010: color_data = 12'b111011101110;
20'b00101100100111011011: color_data = 12'b111011101110;
20'b00101100100111011100: color_data = 12'b111011101110;
20'b00101100100111011101: color_data = 12'b111011101110;
20'b00101100100111011110: color_data = 12'b111011101110;
20'b00101100100111100000: color_data = 12'b111011101110;
20'b00101100100111100001: color_data = 12'b111011101110;
20'b00101100100111100010: color_data = 12'b111011101110;
20'b00101100100111100011: color_data = 12'b111011101110;
20'b00101100100111100100: color_data = 12'b111011101110;
20'b00101100100111100101: color_data = 12'b111011101110;
20'b00101100100111100110: color_data = 12'b111011101110;
20'b00101100100111100111: color_data = 12'b111011101110;
20'b00101100100111101000: color_data = 12'b111011101110;
20'b00101100100111101001: color_data = 12'b111011101110;
20'b00101100110010010110: color_data = 12'b111011101110;
20'b00101100110010010111: color_data = 12'b111011101110;
20'b00101100110010011000: color_data = 12'b111011101110;
20'b00101100110010011001: color_data = 12'b111011101110;
20'b00101100110010011010: color_data = 12'b111011101110;
20'b00101100110010011011: color_data = 12'b111011101110;
20'b00101100110010011100: color_data = 12'b111011101110;
20'b00101100110010011101: color_data = 12'b111011101110;
20'b00101100110010011110: color_data = 12'b111011101110;
20'b00101100110010011111: color_data = 12'b111011101110;
20'b00101100110010100001: color_data = 12'b111011101110;
20'b00101100110010100010: color_data = 12'b111011101110;
20'b00101100110010100011: color_data = 12'b111011101110;
20'b00101100110010100100: color_data = 12'b111011101110;
20'b00101100110010100101: color_data = 12'b111011101110;
20'b00101100110010100110: color_data = 12'b111011101110;
20'b00101100110010100111: color_data = 12'b111011101110;
20'b00101100110010101000: color_data = 12'b111011101110;
20'b00101100110010101001: color_data = 12'b111011101110;
20'b00101100110010101010: color_data = 12'b111011101110;
20'b00101100110010101100: color_data = 12'b111011101110;
20'b00101100110010101101: color_data = 12'b111011101110;
20'b00101100110010101110: color_data = 12'b111011101110;
20'b00101100110010101111: color_data = 12'b111011101110;
20'b00101100110010110000: color_data = 12'b111011101110;
20'b00101100110010110001: color_data = 12'b111011101110;
20'b00101100110010110010: color_data = 12'b111011101110;
20'b00101100110010110011: color_data = 12'b111011101110;
20'b00101100110010110100: color_data = 12'b111011101110;
20'b00101100110010110101: color_data = 12'b111011101110;
20'b00101100110010110111: color_data = 12'b111011101110;
20'b00101100110010111000: color_data = 12'b111011101110;
20'b00101100110010111001: color_data = 12'b111011101110;
20'b00101100110010111010: color_data = 12'b111011101110;
20'b00101100110010111011: color_data = 12'b111011101110;
20'b00101100110010111100: color_data = 12'b111011101110;
20'b00101100110010111101: color_data = 12'b111011101110;
20'b00101100110010111110: color_data = 12'b111011101110;
20'b00101100110010111111: color_data = 12'b111011101110;
20'b00101100110011000000: color_data = 12'b111011101110;
20'b00101100110011000010: color_data = 12'b111011101110;
20'b00101100110011000011: color_data = 12'b111011101110;
20'b00101100110011000100: color_data = 12'b111011101110;
20'b00101100110011000101: color_data = 12'b111011101110;
20'b00101100110011000110: color_data = 12'b111011101110;
20'b00101100110011000111: color_data = 12'b111011101110;
20'b00101100110011001000: color_data = 12'b111011101110;
20'b00101100110011001001: color_data = 12'b111011101110;
20'b00101100110011001010: color_data = 12'b111011101110;
20'b00101100110011001011: color_data = 12'b111011101110;
20'b00101100110011001101: color_data = 12'b111011101110;
20'b00101100110011001110: color_data = 12'b111011101110;
20'b00101100110011001111: color_data = 12'b111011101110;
20'b00101100110011010000: color_data = 12'b111011101110;
20'b00101100110011010001: color_data = 12'b111011101110;
20'b00101100110011010010: color_data = 12'b111011101110;
20'b00101100110011010011: color_data = 12'b111011101110;
20'b00101100110011010100: color_data = 12'b111011101110;
20'b00101100110011010101: color_data = 12'b111011101110;
20'b00101100110011010110: color_data = 12'b111011101110;
20'b00101100110011011000: color_data = 12'b111011101110;
20'b00101100110011011001: color_data = 12'b111011101110;
20'b00101100110011011010: color_data = 12'b111011101110;
20'b00101100110011011011: color_data = 12'b111011101110;
20'b00101100110011011100: color_data = 12'b111011101110;
20'b00101100110011011101: color_data = 12'b111011101110;
20'b00101100110011011110: color_data = 12'b111011101110;
20'b00101100110011011111: color_data = 12'b111011101110;
20'b00101100110011100000: color_data = 12'b111011101110;
20'b00101100110011100001: color_data = 12'b111011101110;
20'b00101100110011101110: color_data = 12'b111011101110;
20'b00101100110011101111: color_data = 12'b111011101110;
20'b00101100110011110000: color_data = 12'b111011101110;
20'b00101100110011110001: color_data = 12'b111011101110;
20'b00101100110011110010: color_data = 12'b111011101110;
20'b00101100110011110011: color_data = 12'b111011101110;
20'b00101100110011110100: color_data = 12'b111011101110;
20'b00101100110011110101: color_data = 12'b111011101110;
20'b00101100110011110110: color_data = 12'b111011101110;
20'b00101100110011110111: color_data = 12'b111011101110;
20'b00101100110011111001: color_data = 12'b111011101110;
20'b00101100110011111010: color_data = 12'b111011101110;
20'b00101100110011111011: color_data = 12'b111011101110;
20'b00101100110011111100: color_data = 12'b111011101110;
20'b00101100110011111101: color_data = 12'b111011101110;
20'b00101100110011111110: color_data = 12'b111011101110;
20'b00101100110011111111: color_data = 12'b111011101110;
20'b00101100110100000000: color_data = 12'b111011101110;
20'b00101100110100000001: color_data = 12'b111011101110;
20'b00101100110100000010: color_data = 12'b111011101110;
20'b00101100110100100101: color_data = 12'b111011101110;
20'b00101100110100100110: color_data = 12'b111011101110;
20'b00101100110100100111: color_data = 12'b111011101110;
20'b00101100110100101000: color_data = 12'b111011101110;
20'b00101100110100101001: color_data = 12'b111011101110;
20'b00101100110100101010: color_data = 12'b111011101110;
20'b00101100110100101011: color_data = 12'b111011101110;
20'b00101100110100101100: color_data = 12'b111011101110;
20'b00101100110100101101: color_data = 12'b111011101110;
20'b00101100110100101110: color_data = 12'b111011101110;
20'b00101100110100110000: color_data = 12'b111011101110;
20'b00101100110100110001: color_data = 12'b111011101110;
20'b00101100110100110010: color_data = 12'b111011101110;
20'b00101100110100110011: color_data = 12'b111011101110;
20'b00101100110100110100: color_data = 12'b111011101110;
20'b00101100110100110101: color_data = 12'b111011101110;
20'b00101100110100110110: color_data = 12'b111011101110;
20'b00101100110100110111: color_data = 12'b111011101110;
20'b00101100110100111000: color_data = 12'b111011101110;
20'b00101100110100111001: color_data = 12'b111011101110;
20'b00101100110101000110: color_data = 12'b111011101110;
20'b00101100110101000111: color_data = 12'b111011101110;
20'b00101100110101001000: color_data = 12'b111011101110;
20'b00101100110101001001: color_data = 12'b111011101110;
20'b00101100110101001010: color_data = 12'b111011101110;
20'b00101100110101001011: color_data = 12'b111011101110;
20'b00101100110101001100: color_data = 12'b111011101110;
20'b00101100110101001101: color_data = 12'b111011101110;
20'b00101100110101001110: color_data = 12'b111011101110;
20'b00101100110101001111: color_data = 12'b111011101110;
20'b00101100110101010001: color_data = 12'b111011101110;
20'b00101100110101010010: color_data = 12'b111011101110;
20'b00101100110101010011: color_data = 12'b111011101110;
20'b00101100110101010100: color_data = 12'b111011101110;
20'b00101100110101010101: color_data = 12'b111011101110;
20'b00101100110101010110: color_data = 12'b111011101110;
20'b00101100110101010111: color_data = 12'b111011101110;
20'b00101100110101011000: color_data = 12'b111011101110;
20'b00101100110101011001: color_data = 12'b111011101110;
20'b00101100110101011010: color_data = 12'b111011101110;
20'b00101100110101111101: color_data = 12'b111011101110;
20'b00101100110101111110: color_data = 12'b111011101110;
20'b00101100110101111111: color_data = 12'b111011101110;
20'b00101100110110000000: color_data = 12'b111011101110;
20'b00101100110110000001: color_data = 12'b111011101110;
20'b00101100110110000010: color_data = 12'b111011101110;
20'b00101100110110000011: color_data = 12'b111011101110;
20'b00101100110110000100: color_data = 12'b111011101110;
20'b00101100110110000101: color_data = 12'b111011101110;
20'b00101100110110000110: color_data = 12'b111011101110;
20'b00101100110110001000: color_data = 12'b111011101110;
20'b00101100110110001001: color_data = 12'b111011101110;
20'b00101100110110001010: color_data = 12'b111011101110;
20'b00101100110110001011: color_data = 12'b111011101110;
20'b00101100110110001100: color_data = 12'b111011101110;
20'b00101100110110001101: color_data = 12'b111011101110;
20'b00101100110110001110: color_data = 12'b111011101110;
20'b00101100110110001111: color_data = 12'b111011101110;
20'b00101100110110010000: color_data = 12'b111011101110;
20'b00101100110110010001: color_data = 12'b111011101110;
20'b00101100110110011110: color_data = 12'b111011101110;
20'b00101100110110011111: color_data = 12'b111011101110;
20'b00101100110110100000: color_data = 12'b111011101110;
20'b00101100110110100001: color_data = 12'b111011101110;
20'b00101100110110100010: color_data = 12'b111011101110;
20'b00101100110110100011: color_data = 12'b111011101110;
20'b00101100110110100100: color_data = 12'b111011101110;
20'b00101100110110100101: color_data = 12'b111011101110;
20'b00101100110110100110: color_data = 12'b111011101110;
20'b00101100110110100111: color_data = 12'b111011101110;
20'b00101100110110101001: color_data = 12'b111011101110;
20'b00101100110110101010: color_data = 12'b111011101110;
20'b00101100110110101011: color_data = 12'b111011101110;
20'b00101100110110101100: color_data = 12'b111011101110;
20'b00101100110110101101: color_data = 12'b111011101110;
20'b00101100110110101110: color_data = 12'b111011101110;
20'b00101100110110101111: color_data = 12'b111011101110;
20'b00101100110110110000: color_data = 12'b111011101110;
20'b00101100110110110001: color_data = 12'b111011101110;
20'b00101100110110110010: color_data = 12'b111011101110;
20'b00101100110110110100: color_data = 12'b111011101110;
20'b00101100110110110101: color_data = 12'b111011101110;
20'b00101100110110110110: color_data = 12'b111011101110;
20'b00101100110110110111: color_data = 12'b111011101110;
20'b00101100110110111000: color_data = 12'b111011101110;
20'b00101100110110111001: color_data = 12'b111011101110;
20'b00101100110110111010: color_data = 12'b111011101110;
20'b00101100110110111011: color_data = 12'b111011101110;
20'b00101100110110111100: color_data = 12'b111011101110;
20'b00101100110110111101: color_data = 12'b111011101110;
20'b00101100110110111111: color_data = 12'b111011101110;
20'b00101100110111000000: color_data = 12'b111011101110;
20'b00101100110111000001: color_data = 12'b111011101110;
20'b00101100110111000010: color_data = 12'b111011101110;
20'b00101100110111000011: color_data = 12'b111011101110;
20'b00101100110111000100: color_data = 12'b111011101110;
20'b00101100110111000101: color_data = 12'b111011101110;
20'b00101100110111000110: color_data = 12'b111011101110;
20'b00101100110111000111: color_data = 12'b111011101110;
20'b00101100110111001000: color_data = 12'b111011101110;
20'b00101100110111001010: color_data = 12'b111011101110;
20'b00101100110111001011: color_data = 12'b111011101110;
20'b00101100110111001100: color_data = 12'b111011101110;
20'b00101100110111001101: color_data = 12'b111011101110;
20'b00101100110111001110: color_data = 12'b111011101110;
20'b00101100110111001111: color_data = 12'b111011101110;
20'b00101100110111010000: color_data = 12'b111011101110;
20'b00101100110111010001: color_data = 12'b111011101110;
20'b00101100110111010010: color_data = 12'b111011101110;
20'b00101100110111010011: color_data = 12'b111011101110;
20'b00101100110111010101: color_data = 12'b111011101110;
20'b00101100110111010110: color_data = 12'b111011101110;
20'b00101100110111010111: color_data = 12'b111011101110;
20'b00101100110111011000: color_data = 12'b111011101110;
20'b00101100110111011001: color_data = 12'b111011101110;
20'b00101100110111011010: color_data = 12'b111011101110;
20'b00101100110111011011: color_data = 12'b111011101110;
20'b00101100110111011100: color_data = 12'b111011101110;
20'b00101100110111011101: color_data = 12'b111011101110;
20'b00101100110111011110: color_data = 12'b111011101110;
20'b00101100110111100000: color_data = 12'b111011101110;
20'b00101100110111100001: color_data = 12'b111011101110;
20'b00101100110111100010: color_data = 12'b111011101110;
20'b00101100110111100011: color_data = 12'b111011101110;
20'b00101100110111100100: color_data = 12'b111011101110;
20'b00101100110111100101: color_data = 12'b111011101110;
20'b00101100110111100110: color_data = 12'b111011101110;
20'b00101100110111100111: color_data = 12'b111011101110;
20'b00101100110111101000: color_data = 12'b111011101110;
20'b00101100110111101001: color_data = 12'b111011101110;
20'b00101101000010010110: color_data = 12'b111011101110;
20'b00101101000010010111: color_data = 12'b111011101110;
20'b00101101000010011000: color_data = 12'b111011101110;
20'b00101101000010011001: color_data = 12'b111011101110;
20'b00101101000010011010: color_data = 12'b111011101110;
20'b00101101000010011011: color_data = 12'b111011101110;
20'b00101101000010011100: color_data = 12'b111011101110;
20'b00101101000010011101: color_data = 12'b111011101110;
20'b00101101000010011110: color_data = 12'b111011101110;
20'b00101101000010011111: color_data = 12'b111011101110;
20'b00101101000010100001: color_data = 12'b111011101110;
20'b00101101000010100010: color_data = 12'b111011101110;
20'b00101101000010100011: color_data = 12'b111011101110;
20'b00101101000010100100: color_data = 12'b111011101110;
20'b00101101000010100101: color_data = 12'b111011101110;
20'b00101101000010100110: color_data = 12'b111011101110;
20'b00101101000010100111: color_data = 12'b111011101110;
20'b00101101000010101000: color_data = 12'b111011101110;
20'b00101101000010101001: color_data = 12'b111011101110;
20'b00101101000010101010: color_data = 12'b111011101110;
20'b00101101000010101100: color_data = 12'b111011101110;
20'b00101101000010101101: color_data = 12'b111011101110;
20'b00101101000010101110: color_data = 12'b111011101110;
20'b00101101000010101111: color_data = 12'b111011101110;
20'b00101101000010110000: color_data = 12'b111011101110;
20'b00101101000010110001: color_data = 12'b111011101110;
20'b00101101000010110010: color_data = 12'b111011101110;
20'b00101101000010110011: color_data = 12'b111011101110;
20'b00101101000010110100: color_data = 12'b111011101110;
20'b00101101000010110101: color_data = 12'b111011101110;
20'b00101101000010110111: color_data = 12'b111011101110;
20'b00101101000010111000: color_data = 12'b111011101110;
20'b00101101000010111001: color_data = 12'b111011101110;
20'b00101101000010111010: color_data = 12'b111011101110;
20'b00101101000010111011: color_data = 12'b111011101110;
20'b00101101000010111100: color_data = 12'b111011101110;
20'b00101101000010111101: color_data = 12'b111011101110;
20'b00101101000010111110: color_data = 12'b111011101110;
20'b00101101000010111111: color_data = 12'b111011101110;
20'b00101101000011000000: color_data = 12'b111011101110;
20'b00101101000011000010: color_data = 12'b111011101110;
20'b00101101000011000011: color_data = 12'b111011101110;
20'b00101101000011000100: color_data = 12'b111011101110;
20'b00101101000011000101: color_data = 12'b111011101110;
20'b00101101000011000110: color_data = 12'b111011101110;
20'b00101101000011000111: color_data = 12'b111011101110;
20'b00101101000011001000: color_data = 12'b111011101110;
20'b00101101000011001001: color_data = 12'b111011101110;
20'b00101101000011001010: color_data = 12'b111011101110;
20'b00101101000011001011: color_data = 12'b111011101110;
20'b00101101000011001101: color_data = 12'b111011101110;
20'b00101101000011001110: color_data = 12'b111011101110;
20'b00101101000011001111: color_data = 12'b111011101110;
20'b00101101000011010000: color_data = 12'b111011101110;
20'b00101101000011010001: color_data = 12'b111011101110;
20'b00101101000011010010: color_data = 12'b111011101110;
20'b00101101000011010011: color_data = 12'b111011101110;
20'b00101101000011010100: color_data = 12'b111011101110;
20'b00101101000011010101: color_data = 12'b111011101110;
20'b00101101000011010110: color_data = 12'b111011101110;
20'b00101101000011011000: color_data = 12'b111011101110;
20'b00101101000011011001: color_data = 12'b111011101110;
20'b00101101000011011010: color_data = 12'b111011101110;
20'b00101101000011011011: color_data = 12'b111011101110;
20'b00101101000011011100: color_data = 12'b111011101110;
20'b00101101000011011101: color_data = 12'b111011101110;
20'b00101101000011011110: color_data = 12'b111011101110;
20'b00101101000011011111: color_data = 12'b111011101110;
20'b00101101000011100000: color_data = 12'b111011101110;
20'b00101101000011100001: color_data = 12'b111011101110;
20'b00101101000011101110: color_data = 12'b111011101110;
20'b00101101000011101111: color_data = 12'b111011101110;
20'b00101101000011110000: color_data = 12'b111011101110;
20'b00101101000011110001: color_data = 12'b111011101110;
20'b00101101000011110010: color_data = 12'b111011101110;
20'b00101101000011110011: color_data = 12'b111011101110;
20'b00101101000011110100: color_data = 12'b111011101110;
20'b00101101000011110101: color_data = 12'b111011101110;
20'b00101101000011110110: color_data = 12'b111011101110;
20'b00101101000011110111: color_data = 12'b111011101110;
20'b00101101000011111001: color_data = 12'b111011101110;
20'b00101101000011111010: color_data = 12'b111011101110;
20'b00101101000011111011: color_data = 12'b111011101110;
20'b00101101000011111100: color_data = 12'b111011101110;
20'b00101101000011111101: color_data = 12'b111011101110;
20'b00101101000011111110: color_data = 12'b111011101110;
20'b00101101000011111111: color_data = 12'b111011101110;
20'b00101101000100000000: color_data = 12'b111011101110;
20'b00101101000100000001: color_data = 12'b111011101110;
20'b00101101000100000010: color_data = 12'b111011101110;
20'b00101101000100100101: color_data = 12'b111011101110;
20'b00101101000100100110: color_data = 12'b111011101110;
20'b00101101000100100111: color_data = 12'b111011101110;
20'b00101101000100101000: color_data = 12'b111011101110;
20'b00101101000100101001: color_data = 12'b111011101110;
20'b00101101000100101010: color_data = 12'b111011101110;
20'b00101101000100101011: color_data = 12'b111011101110;
20'b00101101000100101100: color_data = 12'b111011101110;
20'b00101101000100101101: color_data = 12'b111011101110;
20'b00101101000100101110: color_data = 12'b111011101110;
20'b00101101000100110000: color_data = 12'b111011101110;
20'b00101101000100110001: color_data = 12'b111011101110;
20'b00101101000100110010: color_data = 12'b111011101110;
20'b00101101000100110011: color_data = 12'b111011101110;
20'b00101101000100110100: color_data = 12'b111011101110;
20'b00101101000100110101: color_data = 12'b111011101110;
20'b00101101000100110110: color_data = 12'b111011101110;
20'b00101101000100110111: color_data = 12'b111011101110;
20'b00101101000100111000: color_data = 12'b111011101110;
20'b00101101000100111001: color_data = 12'b111011101110;
20'b00101101000101000110: color_data = 12'b111011101110;
20'b00101101000101000111: color_data = 12'b111011101110;
20'b00101101000101001000: color_data = 12'b111011101110;
20'b00101101000101001001: color_data = 12'b111011101110;
20'b00101101000101001010: color_data = 12'b111011101110;
20'b00101101000101001011: color_data = 12'b111011101110;
20'b00101101000101001100: color_data = 12'b111011101110;
20'b00101101000101001101: color_data = 12'b111011101110;
20'b00101101000101001110: color_data = 12'b111011101110;
20'b00101101000101001111: color_data = 12'b111011101110;
20'b00101101000101010001: color_data = 12'b111011101110;
20'b00101101000101010010: color_data = 12'b111011101110;
20'b00101101000101010011: color_data = 12'b111011101110;
20'b00101101000101010100: color_data = 12'b111011101110;
20'b00101101000101010101: color_data = 12'b111011101110;
20'b00101101000101010110: color_data = 12'b111011101110;
20'b00101101000101010111: color_data = 12'b111011101110;
20'b00101101000101011000: color_data = 12'b111011101110;
20'b00101101000101011001: color_data = 12'b111011101110;
20'b00101101000101011010: color_data = 12'b111011101110;
20'b00101101000101111101: color_data = 12'b111011101110;
20'b00101101000101111110: color_data = 12'b111011101110;
20'b00101101000101111111: color_data = 12'b111011101110;
20'b00101101000110000000: color_data = 12'b111011101110;
20'b00101101000110000001: color_data = 12'b111011101110;
20'b00101101000110000010: color_data = 12'b111011101110;
20'b00101101000110000011: color_data = 12'b111011101110;
20'b00101101000110000100: color_data = 12'b111011101110;
20'b00101101000110000101: color_data = 12'b111011101110;
20'b00101101000110000110: color_data = 12'b111011101110;
20'b00101101000110001000: color_data = 12'b111011101110;
20'b00101101000110001001: color_data = 12'b111011101110;
20'b00101101000110001010: color_data = 12'b111011101110;
20'b00101101000110001011: color_data = 12'b111011101110;
20'b00101101000110001100: color_data = 12'b111011101110;
20'b00101101000110001101: color_data = 12'b111011101110;
20'b00101101000110001110: color_data = 12'b111011101110;
20'b00101101000110001111: color_data = 12'b111011101110;
20'b00101101000110010000: color_data = 12'b111011101110;
20'b00101101000110010001: color_data = 12'b111011101110;
20'b00101101000110011110: color_data = 12'b111011101110;
20'b00101101000110011111: color_data = 12'b111011101110;
20'b00101101000110100000: color_data = 12'b111011101110;
20'b00101101000110100001: color_data = 12'b111011101110;
20'b00101101000110100010: color_data = 12'b111011101110;
20'b00101101000110100011: color_data = 12'b111011101110;
20'b00101101000110100100: color_data = 12'b111011101110;
20'b00101101000110100101: color_data = 12'b111011101110;
20'b00101101000110100110: color_data = 12'b111011101110;
20'b00101101000110100111: color_data = 12'b111011101110;
20'b00101101000110101001: color_data = 12'b111011101110;
20'b00101101000110101010: color_data = 12'b111011101110;
20'b00101101000110101011: color_data = 12'b111011101110;
20'b00101101000110101100: color_data = 12'b111011101110;
20'b00101101000110101101: color_data = 12'b111011101110;
20'b00101101000110101110: color_data = 12'b111011101110;
20'b00101101000110101111: color_data = 12'b111011101110;
20'b00101101000110110000: color_data = 12'b111011101110;
20'b00101101000110110001: color_data = 12'b111011101110;
20'b00101101000110110010: color_data = 12'b111011101110;
20'b00101101000110110100: color_data = 12'b111011101110;
20'b00101101000110110101: color_data = 12'b111011101110;
20'b00101101000110110110: color_data = 12'b111011101110;
20'b00101101000110110111: color_data = 12'b111011101110;
20'b00101101000110111000: color_data = 12'b111011101110;
20'b00101101000110111001: color_data = 12'b111011101110;
20'b00101101000110111010: color_data = 12'b111011101110;
20'b00101101000110111011: color_data = 12'b111011101110;
20'b00101101000110111100: color_data = 12'b111011101110;
20'b00101101000110111101: color_data = 12'b111011101110;
20'b00101101000110111111: color_data = 12'b111011101110;
20'b00101101000111000000: color_data = 12'b111011101110;
20'b00101101000111000001: color_data = 12'b111011101110;
20'b00101101000111000010: color_data = 12'b111011101110;
20'b00101101000111000011: color_data = 12'b111011101110;
20'b00101101000111000100: color_data = 12'b111011101110;
20'b00101101000111000101: color_data = 12'b111011101110;
20'b00101101000111000110: color_data = 12'b111011101110;
20'b00101101000111000111: color_data = 12'b111011101110;
20'b00101101000111001000: color_data = 12'b111011101110;
20'b00101101000111001010: color_data = 12'b111011101110;
20'b00101101000111001011: color_data = 12'b111011101110;
20'b00101101000111001100: color_data = 12'b111011101110;
20'b00101101000111001101: color_data = 12'b111011101110;
20'b00101101000111001110: color_data = 12'b111011101110;
20'b00101101000111001111: color_data = 12'b111011101110;
20'b00101101000111010000: color_data = 12'b111011101110;
20'b00101101000111010001: color_data = 12'b111011101110;
20'b00101101000111010010: color_data = 12'b111011101110;
20'b00101101000111010011: color_data = 12'b111011101110;
20'b00101101000111010101: color_data = 12'b111011101110;
20'b00101101000111010110: color_data = 12'b111011101110;
20'b00101101000111010111: color_data = 12'b111011101110;
20'b00101101000111011000: color_data = 12'b111011101110;
20'b00101101000111011001: color_data = 12'b111011101110;
20'b00101101000111011010: color_data = 12'b111011101110;
20'b00101101000111011011: color_data = 12'b111011101110;
20'b00101101000111011100: color_data = 12'b111011101110;
20'b00101101000111011101: color_data = 12'b111011101110;
20'b00101101000111011110: color_data = 12'b111011101110;
20'b00101101000111100000: color_data = 12'b111011101110;
20'b00101101000111100001: color_data = 12'b111011101110;
20'b00101101000111100010: color_data = 12'b111011101110;
20'b00101101000111100011: color_data = 12'b111011101110;
20'b00101101000111100100: color_data = 12'b111011101110;
20'b00101101000111100101: color_data = 12'b111011101110;
20'b00101101000111100110: color_data = 12'b111011101110;
20'b00101101000111100111: color_data = 12'b111011101110;
20'b00101101000111101000: color_data = 12'b111011101110;
20'b00101101000111101001: color_data = 12'b111011101110;
20'b00101101010010010110: color_data = 12'b111011101110;
20'b00101101010010010111: color_data = 12'b111011101110;
20'b00101101010010011000: color_data = 12'b111011101110;
20'b00101101010010011001: color_data = 12'b111011101110;
20'b00101101010010011010: color_data = 12'b111011101110;
20'b00101101010010011011: color_data = 12'b111011101110;
20'b00101101010010011100: color_data = 12'b111011101110;
20'b00101101010010011101: color_data = 12'b111011101110;
20'b00101101010010011110: color_data = 12'b111011101110;
20'b00101101010010011111: color_data = 12'b111011101110;
20'b00101101010010100001: color_data = 12'b111011101110;
20'b00101101010010100010: color_data = 12'b111011101110;
20'b00101101010010100011: color_data = 12'b111011101110;
20'b00101101010010100100: color_data = 12'b111011101110;
20'b00101101010010100101: color_data = 12'b111011101110;
20'b00101101010010100110: color_data = 12'b111011101110;
20'b00101101010010100111: color_data = 12'b111011101110;
20'b00101101010010101000: color_data = 12'b111011101110;
20'b00101101010010101001: color_data = 12'b111011101110;
20'b00101101010010101010: color_data = 12'b111011101110;
20'b00101101010010101100: color_data = 12'b111011101110;
20'b00101101010010101101: color_data = 12'b111011101110;
20'b00101101010010101110: color_data = 12'b111011101110;
20'b00101101010010101111: color_data = 12'b111011101110;
20'b00101101010010110000: color_data = 12'b111011101110;
20'b00101101010010110001: color_data = 12'b111011101110;
20'b00101101010010110010: color_data = 12'b111011101110;
20'b00101101010010110011: color_data = 12'b111011101110;
20'b00101101010010110100: color_data = 12'b111011101110;
20'b00101101010010110101: color_data = 12'b111011101110;
20'b00101101010010110111: color_data = 12'b111011101110;
20'b00101101010010111000: color_data = 12'b111011101110;
20'b00101101010010111001: color_data = 12'b111011101110;
20'b00101101010010111010: color_data = 12'b111011101110;
20'b00101101010010111011: color_data = 12'b111011101110;
20'b00101101010010111100: color_data = 12'b111011101110;
20'b00101101010010111101: color_data = 12'b111011101110;
20'b00101101010010111110: color_data = 12'b111011101110;
20'b00101101010010111111: color_data = 12'b111011101110;
20'b00101101010011000000: color_data = 12'b111011101110;
20'b00101101010011000010: color_data = 12'b111011101110;
20'b00101101010011000011: color_data = 12'b111011101110;
20'b00101101010011000100: color_data = 12'b111011101110;
20'b00101101010011000101: color_data = 12'b111011101110;
20'b00101101010011000110: color_data = 12'b111011101110;
20'b00101101010011000111: color_data = 12'b111011101110;
20'b00101101010011001000: color_data = 12'b111011101110;
20'b00101101010011001001: color_data = 12'b111011101110;
20'b00101101010011001010: color_data = 12'b111011101110;
20'b00101101010011001011: color_data = 12'b111011101110;
20'b00101101010011001101: color_data = 12'b111011101110;
20'b00101101010011001110: color_data = 12'b111011101110;
20'b00101101010011001111: color_data = 12'b111011101110;
20'b00101101010011010000: color_data = 12'b111011101110;
20'b00101101010011010001: color_data = 12'b111011101110;
20'b00101101010011010010: color_data = 12'b111011101110;
20'b00101101010011010011: color_data = 12'b111011101110;
20'b00101101010011010100: color_data = 12'b111011101110;
20'b00101101010011010101: color_data = 12'b111011101110;
20'b00101101010011010110: color_data = 12'b111011101110;
20'b00101101010011011000: color_data = 12'b111011101110;
20'b00101101010011011001: color_data = 12'b111011101110;
20'b00101101010011011010: color_data = 12'b111011101110;
20'b00101101010011011011: color_data = 12'b111011101110;
20'b00101101010011011100: color_data = 12'b111011101110;
20'b00101101010011011101: color_data = 12'b111011101110;
20'b00101101010011011110: color_data = 12'b111011101110;
20'b00101101010011011111: color_data = 12'b111011101110;
20'b00101101010011100000: color_data = 12'b111011101110;
20'b00101101010011100001: color_data = 12'b111011101110;
20'b00101101010011101110: color_data = 12'b111011101110;
20'b00101101010011101111: color_data = 12'b111011101110;
20'b00101101010011110000: color_data = 12'b111011101110;
20'b00101101010011110001: color_data = 12'b111011101110;
20'b00101101010011110010: color_data = 12'b111011101110;
20'b00101101010011110011: color_data = 12'b111011101110;
20'b00101101010011110100: color_data = 12'b111011101110;
20'b00101101010011110101: color_data = 12'b111011101110;
20'b00101101010011110110: color_data = 12'b111011101110;
20'b00101101010011110111: color_data = 12'b111011101110;
20'b00101101010011111001: color_data = 12'b111011101110;
20'b00101101010011111010: color_data = 12'b111011101110;
20'b00101101010011111011: color_data = 12'b111011101110;
20'b00101101010011111100: color_data = 12'b111011101110;
20'b00101101010011111101: color_data = 12'b111011101110;
20'b00101101010011111110: color_data = 12'b111011101110;
20'b00101101010011111111: color_data = 12'b111011101110;
20'b00101101010100000000: color_data = 12'b111011101110;
20'b00101101010100000001: color_data = 12'b111011101110;
20'b00101101010100000010: color_data = 12'b111011101110;
20'b00101101010100100101: color_data = 12'b111011101110;
20'b00101101010100100110: color_data = 12'b111011101110;
20'b00101101010100100111: color_data = 12'b111011101110;
20'b00101101010100101000: color_data = 12'b111011101110;
20'b00101101010100101001: color_data = 12'b111011101110;
20'b00101101010100101010: color_data = 12'b111011101110;
20'b00101101010100101011: color_data = 12'b111011101110;
20'b00101101010100101100: color_data = 12'b111011101110;
20'b00101101010100101101: color_data = 12'b111011101110;
20'b00101101010100101110: color_data = 12'b111011101110;
20'b00101101010100110000: color_data = 12'b111011101110;
20'b00101101010100110001: color_data = 12'b111011101110;
20'b00101101010100110010: color_data = 12'b111011101110;
20'b00101101010100110011: color_data = 12'b111011101110;
20'b00101101010100110100: color_data = 12'b111011101110;
20'b00101101010100110101: color_data = 12'b111011101110;
20'b00101101010100110110: color_data = 12'b111011101110;
20'b00101101010100110111: color_data = 12'b111011101110;
20'b00101101010100111000: color_data = 12'b111011101110;
20'b00101101010100111001: color_data = 12'b111011101110;
20'b00101101010101000110: color_data = 12'b111011101110;
20'b00101101010101000111: color_data = 12'b111011101110;
20'b00101101010101001000: color_data = 12'b111011101110;
20'b00101101010101001001: color_data = 12'b111011101110;
20'b00101101010101001010: color_data = 12'b111011101110;
20'b00101101010101001011: color_data = 12'b111011101110;
20'b00101101010101001100: color_data = 12'b111011101110;
20'b00101101010101001101: color_data = 12'b111011101110;
20'b00101101010101001110: color_data = 12'b111011101110;
20'b00101101010101001111: color_data = 12'b111011101110;
20'b00101101010101010001: color_data = 12'b111011101110;
20'b00101101010101010010: color_data = 12'b111011101110;
20'b00101101010101010011: color_data = 12'b111011101110;
20'b00101101010101010100: color_data = 12'b111011101110;
20'b00101101010101010101: color_data = 12'b111011101110;
20'b00101101010101010110: color_data = 12'b111011101110;
20'b00101101010101010111: color_data = 12'b111011101110;
20'b00101101010101011000: color_data = 12'b111011101110;
20'b00101101010101011001: color_data = 12'b111011101110;
20'b00101101010101011010: color_data = 12'b111011101110;
20'b00101101010101111101: color_data = 12'b111011101110;
20'b00101101010101111110: color_data = 12'b111011101110;
20'b00101101010101111111: color_data = 12'b111011101110;
20'b00101101010110000000: color_data = 12'b111011101110;
20'b00101101010110000001: color_data = 12'b111011101110;
20'b00101101010110000010: color_data = 12'b111011101110;
20'b00101101010110000011: color_data = 12'b111011101110;
20'b00101101010110000100: color_data = 12'b111011101110;
20'b00101101010110000101: color_data = 12'b111011101110;
20'b00101101010110000110: color_data = 12'b111011101110;
20'b00101101010110001000: color_data = 12'b111011101110;
20'b00101101010110001001: color_data = 12'b111011101110;
20'b00101101010110001010: color_data = 12'b111011101110;
20'b00101101010110001011: color_data = 12'b111011101110;
20'b00101101010110001100: color_data = 12'b111011101110;
20'b00101101010110001101: color_data = 12'b111011101110;
20'b00101101010110001110: color_data = 12'b111011101110;
20'b00101101010110001111: color_data = 12'b111011101110;
20'b00101101010110010000: color_data = 12'b111011101110;
20'b00101101010110010001: color_data = 12'b111011101110;
20'b00101101010110011110: color_data = 12'b111011101110;
20'b00101101010110011111: color_data = 12'b111011101110;
20'b00101101010110100000: color_data = 12'b111011101110;
20'b00101101010110100001: color_data = 12'b111011101110;
20'b00101101010110100010: color_data = 12'b111011101110;
20'b00101101010110100011: color_data = 12'b111011101110;
20'b00101101010110100100: color_data = 12'b111011101110;
20'b00101101010110100101: color_data = 12'b111011101110;
20'b00101101010110100110: color_data = 12'b111011101110;
20'b00101101010110100111: color_data = 12'b111011101110;
20'b00101101010110101001: color_data = 12'b111011101110;
20'b00101101010110101010: color_data = 12'b111011101110;
20'b00101101010110101011: color_data = 12'b111011101110;
20'b00101101010110101100: color_data = 12'b111011101110;
20'b00101101010110101101: color_data = 12'b111011101110;
20'b00101101010110101110: color_data = 12'b111011101110;
20'b00101101010110101111: color_data = 12'b111011101110;
20'b00101101010110110000: color_data = 12'b111011101110;
20'b00101101010110110001: color_data = 12'b111011101110;
20'b00101101010110110010: color_data = 12'b111011101110;
20'b00101101010110110100: color_data = 12'b111011101110;
20'b00101101010110110101: color_data = 12'b111011101110;
20'b00101101010110110110: color_data = 12'b111011101110;
20'b00101101010110110111: color_data = 12'b111011101110;
20'b00101101010110111000: color_data = 12'b111011101110;
20'b00101101010110111001: color_data = 12'b111011101110;
20'b00101101010110111010: color_data = 12'b111011101110;
20'b00101101010110111011: color_data = 12'b111011101110;
20'b00101101010110111100: color_data = 12'b111011101110;
20'b00101101010110111101: color_data = 12'b111011101110;
20'b00101101010110111111: color_data = 12'b111011101110;
20'b00101101010111000000: color_data = 12'b111011101110;
20'b00101101010111000001: color_data = 12'b111011101110;
20'b00101101010111000010: color_data = 12'b111011101110;
20'b00101101010111000011: color_data = 12'b111011101110;
20'b00101101010111000100: color_data = 12'b111011101110;
20'b00101101010111000101: color_data = 12'b111011101110;
20'b00101101010111000110: color_data = 12'b111011101110;
20'b00101101010111000111: color_data = 12'b111011101110;
20'b00101101010111001000: color_data = 12'b111011101110;
20'b00101101010111001010: color_data = 12'b111011101110;
20'b00101101010111001011: color_data = 12'b111011101110;
20'b00101101010111001100: color_data = 12'b111011101110;
20'b00101101010111001101: color_data = 12'b111011101110;
20'b00101101010111001110: color_data = 12'b111011101110;
20'b00101101010111001111: color_data = 12'b111011101110;
20'b00101101010111010000: color_data = 12'b111011101110;
20'b00101101010111010001: color_data = 12'b111011101110;
20'b00101101010111010010: color_data = 12'b111011101110;
20'b00101101010111010011: color_data = 12'b111011101110;
20'b00101101010111010101: color_data = 12'b111011101110;
20'b00101101010111010110: color_data = 12'b111011101110;
20'b00101101010111010111: color_data = 12'b111011101110;
20'b00101101010111011000: color_data = 12'b111011101110;
20'b00101101010111011001: color_data = 12'b111011101110;
20'b00101101010111011010: color_data = 12'b111011101110;
20'b00101101010111011011: color_data = 12'b111011101110;
20'b00101101010111011100: color_data = 12'b111011101110;
20'b00101101010111011101: color_data = 12'b111011101110;
20'b00101101010111011110: color_data = 12'b111011101110;
20'b00101101010111100000: color_data = 12'b111011101110;
20'b00101101010111100001: color_data = 12'b111011101110;
20'b00101101010111100010: color_data = 12'b111011101110;
20'b00101101010111100011: color_data = 12'b111011101110;
20'b00101101010111100100: color_data = 12'b111011101110;
20'b00101101010111100101: color_data = 12'b111011101110;
20'b00101101010111100110: color_data = 12'b111011101110;
20'b00101101010111100111: color_data = 12'b111011101110;
20'b00101101010111101000: color_data = 12'b111011101110;
20'b00101101010111101001: color_data = 12'b111011101110;
20'b00101101100010010110: color_data = 12'b111011101110;
20'b00101101100010010111: color_data = 12'b111011101110;
20'b00101101100010011000: color_data = 12'b111011101110;
20'b00101101100010011001: color_data = 12'b111011101110;
20'b00101101100010011010: color_data = 12'b111011101110;
20'b00101101100010011011: color_data = 12'b111011101110;
20'b00101101100010011100: color_data = 12'b111011101110;
20'b00101101100010011101: color_data = 12'b111011101110;
20'b00101101100010011110: color_data = 12'b111011101110;
20'b00101101100010011111: color_data = 12'b111011101110;
20'b00101101100010100001: color_data = 12'b111011101110;
20'b00101101100010100010: color_data = 12'b111011101110;
20'b00101101100010100011: color_data = 12'b111011101110;
20'b00101101100010100100: color_data = 12'b111011101110;
20'b00101101100010100101: color_data = 12'b111011101110;
20'b00101101100010100110: color_data = 12'b111011101110;
20'b00101101100010100111: color_data = 12'b111011101110;
20'b00101101100010101000: color_data = 12'b111011101110;
20'b00101101100010101001: color_data = 12'b111011101110;
20'b00101101100010101010: color_data = 12'b111011101110;
20'b00101101100010101100: color_data = 12'b111011101110;
20'b00101101100010101101: color_data = 12'b111011101110;
20'b00101101100010101110: color_data = 12'b111011101110;
20'b00101101100010101111: color_data = 12'b111011101110;
20'b00101101100010110000: color_data = 12'b111011101110;
20'b00101101100010110001: color_data = 12'b111011101110;
20'b00101101100010110010: color_data = 12'b111011101110;
20'b00101101100010110011: color_data = 12'b111011101110;
20'b00101101100010110100: color_data = 12'b111011101110;
20'b00101101100010110101: color_data = 12'b111011101110;
20'b00101101100010110111: color_data = 12'b111011101110;
20'b00101101100010111000: color_data = 12'b111011101110;
20'b00101101100010111001: color_data = 12'b111011101110;
20'b00101101100010111010: color_data = 12'b111011101110;
20'b00101101100010111011: color_data = 12'b111011101110;
20'b00101101100010111100: color_data = 12'b111011101110;
20'b00101101100010111101: color_data = 12'b111011101110;
20'b00101101100010111110: color_data = 12'b111011101110;
20'b00101101100010111111: color_data = 12'b111011101110;
20'b00101101100011000000: color_data = 12'b111011101110;
20'b00101101100011000010: color_data = 12'b111011101110;
20'b00101101100011000011: color_data = 12'b111011101110;
20'b00101101100011000100: color_data = 12'b111011101110;
20'b00101101100011000101: color_data = 12'b111011101110;
20'b00101101100011000110: color_data = 12'b111011101110;
20'b00101101100011000111: color_data = 12'b111011101110;
20'b00101101100011001000: color_data = 12'b111011101110;
20'b00101101100011001001: color_data = 12'b111011101110;
20'b00101101100011001010: color_data = 12'b111011101110;
20'b00101101100011001011: color_data = 12'b111011101110;
20'b00101101100011001101: color_data = 12'b111011101110;
20'b00101101100011001110: color_data = 12'b111011101110;
20'b00101101100011001111: color_data = 12'b111011101110;
20'b00101101100011010000: color_data = 12'b111011101110;
20'b00101101100011010001: color_data = 12'b111011101110;
20'b00101101100011010010: color_data = 12'b111011101110;
20'b00101101100011010011: color_data = 12'b111011101110;
20'b00101101100011010100: color_data = 12'b111011101110;
20'b00101101100011010101: color_data = 12'b111011101110;
20'b00101101100011010110: color_data = 12'b111011101110;
20'b00101101100011011000: color_data = 12'b111011101110;
20'b00101101100011011001: color_data = 12'b111011101110;
20'b00101101100011011010: color_data = 12'b111011101110;
20'b00101101100011011011: color_data = 12'b111011101110;
20'b00101101100011011100: color_data = 12'b111011101110;
20'b00101101100011011101: color_data = 12'b111011101110;
20'b00101101100011011110: color_data = 12'b111011101110;
20'b00101101100011011111: color_data = 12'b111011101110;
20'b00101101100011100000: color_data = 12'b111011101110;
20'b00101101100011100001: color_data = 12'b111011101110;
20'b00101101100011101110: color_data = 12'b111011101110;
20'b00101101100011101111: color_data = 12'b111011101110;
20'b00101101100011110000: color_data = 12'b111011101110;
20'b00101101100011110001: color_data = 12'b111011101110;
20'b00101101100011110010: color_data = 12'b111011101110;
20'b00101101100011110011: color_data = 12'b111011101110;
20'b00101101100011110100: color_data = 12'b111011101110;
20'b00101101100011110101: color_data = 12'b111011101110;
20'b00101101100011110110: color_data = 12'b111011101110;
20'b00101101100011110111: color_data = 12'b111011101110;
20'b00101101100011111001: color_data = 12'b111011101110;
20'b00101101100011111010: color_data = 12'b111011101110;
20'b00101101100011111011: color_data = 12'b111011101110;
20'b00101101100011111100: color_data = 12'b111011101110;
20'b00101101100011111101: color_data = 12'b111011101110;
20'b00101101100011111110: color_data = 12'b111011101110;
20'b00101101100011111111: color_data = 12'b111011101110;
20'b00101101100100000000: color_data = 12'b111011101110;
20'b00101101100100000001: color_data = 12'b111011101110;
20'b00101101100100000010: color_data = 12'b111011101110;
20'b00101101100100100101: color_data = 12'b111011101110;
20'b00101101100100100110: color_data = 12'b111011101110;
20'b00101101100100100111: color_data = 12'b111011101110;
20'b00101101100100101000: color_data = 12'b111011101110;
20'b00101101100100101001: color_data = 12'b111011101110;
20'b00101101100100101010: color_data = 12'b111011101110;
20'b00101101100100101011: color_data = 12'b111011101110;
20'b00101101100100101100: color_data = 12'b111011101110;
20'b00101101100100101101: color_data = 12'b111011101110;
20'b00101101100100101110: color_data = 12'b111011101110;
20'b00101101100100110000: color_data = 12'b111011101110;
20'b00101101100100110001: color_data = 12'b111011101110;
20'b00101101100100110010: color_data = 12'b111011101110;
20'b00101101100100110011: color_data = 12'b111011101110;
20'b00101101100100110100: color_data = 12'b111011101110;
20'b00101101100100110101: color_data = 12'b111011101110;
20'b00101101100100110110: color_data = 12'b111011101110;
20'b00101101100100110111: color_data = 12'b111011101110;
20'b00101101100100111000: color_data = 12'b111011101110;
20'b00101101100100111001: color_data = 12'b111011101110;
20'b00101101100101000110: color_data = 12'b111011101110;
20'b00101101100101000111: color_data = 12'b111011101110;
20'b00101101100101001000: color_data = 12'b111011101110;
20'b00101101100101001001: color_data = 12'b111011101110;
20'b00101101100101001010: color_data = 12'b111011101110;
20'b00101101100101001011: color_data = 12'b111011101110;
20'b00101101100101001100: color_data = 12'b111011101110;
20'b00101101100101001101: color_data = 12'b111011101110;
20'b00101101100101001110: color_data = 12'b111011101110;
20'b00101101100101001111: color_data = 12'b111011101110;
20'b00101101100101010001: color_data = 12'b111011101110;
20'b00101101100101010010: color_data = 12'b111011101110;
20'b00101101100101010011: color_data = 12'b111011101110;
20'b00101101100101010100: color_data = 12'b111011101110;
20'b00101101100101010101: color_data = 12'b111011101110;
20'b00101101100101010110: color_data = 12'b111011101110;
20'b00101101100101010111: color_data = 12'b111011101110;
20'b00101101100101011000: color_data = 12'b111011101110;
20'b00101101100101011001: color_data = 12'b111011101110;
20'b00101101100101011010: color_data = 12'b111011101110;
20'b00101101100101111101: color_data = 12'b111011101110;
20'b00101101100101111110: color_data = 12'b111011101110;
20'b00101101100101111111: color_data = 12'b111011101110;
20'b00101101100110000000: color_data = 12'b111011101110;
20'b00101101100110000001: color_data = 12'b111011101110;
20'b00101101100110000010: color_data = 12'b111011101110;
20'b00101101100110000011: color_data = 12'b111011101110;
20'b00101101100110000100: color_data = 12'b111011101110;
20'b00101101100110000101: color_data = 12'b111011101110;
20'b00101101100110000110: color_data = 12'b111011101110;
20'b00101101100110001000: color_data = 12'b111011101110;
20'b00101101100110001001: color_data = 12'b111011101110;
20'b00101101100110001010: color_data = 12'b111011101110;
20'b00101101100110001011: color_data = 12'b111011101110;
20'b00101101100110001100: color_data = 12'b111011101110;
20'b00101101100110001101: color_data = 12'b111011101110;
20'b00101101100110001110: color_data = 12'b111011101110;
20'b00101101100110001111: color_data = 12'b111011101110;
20'b00101101100110010000: color_data = 12'b111011101110;
20'b00101101100110010001: color_data = 12'b111011101110;
20'b00101101100110011110: color_data = 12'b111011101110;
20'b00101101100110011111: color_data = 12'b111011101110;
20'b00101101100110100000: color_data = 12'b111011101110;
20'b00101101100110100001: color_data = 12'b111011101110;
20'b00101101100110100010: color_data = 12'b111011101110;
20'b00101101100110100011: color_data = 12'b111011101110;
20'b00101101100110100100: color_data = 12'b111011101110;
20'b00101101100110100101: color_data = 12'b111011101110;
20'b00101101100110100110: color_data = 12'b111011101110;
20'b00101101100110100111: color_data = 12'b111011101110;
20'b00101101100110101001: color_data = 12'b111011101110;
20'b00101101100110101010: color_data = 12'b111011101110;
20'b00101101100110101011: color_data = 12'b111011101110;
20'b00101101100110101100: color_data = 12'b111011101110;
20'b00101101100110101101: color_data = 12'b111011101110;
20'b00101101100110101110: color_data = 12'b111011101110;
20'b00101101100110101111: color_data = 12'b111011101110;
20'b00101101100110110000: color_data = 12'b111011101110;
20'b00101101100110110001: color_data = 12'b111011101110;
20'b00101101100110110010: color_data = 12'b111011101110;
20'b00101101100110110100: color_data = 12'b111011101110;
20'b00101101100110110101: color_data = 12'b111011101110;
20'b00101101100110110110: color_data = 12'b111011101110;
20'b00101101100110110111: color_data = 12'b111011101110;
20'b00101101100110111000: color_data = 12'b111011101110;
20'b00101101100110111001: color_data = 12'b111011101110;
20'b00101101100110111010: color_data = 12'b111011101110;
20'b00101101100110111011: color_data = 12'b111011101110;
20'b00101101100110111100: color_data = 12'b111011101110;
20'b00101101100110111101: color_data = 12'b111011101110;
20'b00101101100110111111: color_data = 12'b111011101110;
20'b00101101100111000000: color_data = 12'b111011101110;
20'b00101101100111000001: color_data = 12'b111011101110;
20'b00101101100111000010: color_data = 12'b111011101110;
20'b00101101100111000011: color_data = 12'b111011101110;
20'b00101101100111000100: color_data = 12'b111011101110;
20'b00101101100111000101: color_data = 12'b111011101110;
20'b00101101100111000110: color_data = 12'b111011101110;
20'b00101101100111000111: color_data = 12'b111011101110;
20'b00101101100111001000: color_data = 12'b111011101110;
20'b00101101100111001010: color_data = 12'b111011101110;
20'b00101101100111001011: color_data = 12'b111011101110;
20'b00101101100111001100: color_data = 12'b111011101110;
20'b00101101100111001101: color_data = 12'b111011101110;
20'b00101101100111001110: color_data = 12'b111011101110;
20'b00101101100111001111: color_data = 12'b111011101110;
20'b00101101100111010000: color_data = 12'b111011101110;
20'b00101101100111010001: color_data = 12'b111011101110;
20'b00101101100111010010: color_data = 12'b111011101110;
20'b00101101100111010011: color_data = 12'b111011101110;
20'b00101101100111010101: color_data = 12'b111011101110;
20'b00101101100111010110: color_data = 12'b111011101110;
20'b00101101100111010111: color_data = 12'b111011101110;
20'b00101101100111011000: color_data = 12'b111011101110;
20'b00101101100111011001: color_data = 12'b111011101110;
20'b00101101100111011010: color_data = 12'b111011101110;
20'b00101101100111011011: color_data = 12'b111011101110;
20'b00101101100111011100: color_data = 12'b111011101110;
20'b00101101100111011101: color_data = 12'b111011101110;
20'b00101101100111011110: color_data = 12'b111011101110;
20'b00101101100111100000: color_data = 12'b111011101110;
20'b00101101100111100001: color_data = 12'b111011101110;
20'b00101101100111100010: color_data = 12'b111011101110;
20'b00101101100111100011: color_data = 12'b111011101110;
20'b00101101100111100100: color_data = 12'b111011101110;
20'b00101101100111100101: color_data = 12'b111011101110;
20'b00101101100111100110: color_data = 12'b111011101110;
20'b00101101100111100111: color_data = 12'b111011101110;
20'b00101101100111101000: color_data = 12'b111011101110;
20'b00101101100111101001: color_data = 12'b111011101110;
20'b00101101110010010110: color_data = 12'b111011101110;
20'b00101101110010010111: color_data = 12'b111011101110;
20'b00101101110010011000: color_data = 12'b111011101110;
20'b00101101110010011001: color_data = 12'b111011101110;
20'b00101101110010011010: color_data = 12'b111011101110;
20'b00101101110010011011: color_data = 12'b111011101110;
20'b00101101110010011100: color_data = 12'b111011101110;
20'b00101101110010011101: color_data = 12'b111011101110;
20'b00101101110010011110: color_data = 12'b111011101110;
20'b00101101110010011111: color_data = 12'b111011101110;
20'b00101101110010100001: color_data = 12'b111011101110;
20'b00101101110010100010: color_data = 12'b111011101110;
20'b00101101110010100011: color_data = 12'b111011101110;
20'b00101101110010100100: color_data = 12'b111011101110;
20'b00101101110010100101: color_data = 12'b111011101110;
20'b00101101110010100110: color_data = 12'b111011101110;
20'b00101101110010100111: color_data = 12'b111011101110;
20'b00101101110010101000: color_data = 12'b111011101110;
20'b00101101110010101001: color_data = 12'b111011101110;
20'b00101101110010101010: color_data = 12'b111011101110;
20'b00101101110010101100: color_data = 12'b111011101110;
20'b00101101110010101101: color_data = 12'b111011101110;
20'b00101101110010101110: color_data = 12'b111011101110;
20'b00101101110010101111: color_data = 12'b111011101110;
20'b00101101110010110000: color_data = 12'b111011101110;
20'b00101101110010110001: color_data = 12'b111011101110;
20'b00101101110010110010: color_data = 12'b111011101110;
20'b00101101110010110011: color_data = 12'b111011101110;
20'b00101101110010110100: color_data = 12'b111011101110;
20'b00101101110010110101: color_data = 12'b111011101110;
20'b00101101110010110111: color_data = 12'b111011101110;
20'b00101101110010111000: color_data = 12'b111011101110;
20'b00101101110010111001: color_data = 12'b111011101110;
20'b00101101110010111010: color_data = 12'b111011101110;
20'b00101101110010111011: color_data = 12'b111011101110;
20'b00101101110010111100: color_data = 12'b111011101110;
20'b00101101110010111101: color_data = 12'b111011101110;
20'b00101101110010111110: color_data = 12'b111011101110;
20'b00101101110010111111: color_data = 12'b111011101110;
20'b00101101110011000000: color_data = 12'b111011101110;
20'b00101101110011000010: color_data = 12'b111011101110;
20'b00101101110011000011: color_data = 12'b111011101110;
20'b00101101110011000100: color_data = 12'b111011101110;
20'b00101101110011000101: color_data = 12'b111011101110;
20'b00101101110011000110: color_data = 12'b111011101110;
20'b00101101110011000111: color_data = 12'b111011101110;
20'b00101101110011001000: color_data = 12'b111011101110;
20'b00101101110011001001: color_data = 12'b111011101110;
20'b00101101110011001010: color_data = 12'b111011101110;
20'b00101101110011001011: color_data = 12'b111011101110;
20'b00101101110011001101: color_data = 12'b111011101110;
20'b00101101110011001110: color_data = 12'b111011101110;
20'b00101101110011001111: color_data = 12'b111011101110;
20'b00101101110011010000: color_data = 12'b111011101110;
20'b00101101110011010001: color_data = 12'b111011101110;
20'b00101101110011010010: color_data = 12'b111011101110;
20'b00101101110011010011: color_data = 12'b111011101110;
20'b00101101110011010100: color_data = 12'b111011101110;
20'b00101101110011010101: color_data = 12'b111011101110;
20'b00101101110011010110: color_data = 12'b111011101110;
20'b00101101110011011000: color_data = 12'b111011101110;
20'b00101101110011011001: color_data = 12'b111011101110;
20'b00101101110011011010: color_data = 12'b111011101110;
20'b00101101110011011011: color_data = 12'b111011101110;
20'b00101101110011011100: color_data = 12'b111011101110;
20'b00101101110011011101: color_data = 12'b111011101110;
20'b00101101110011011110: color_data = 12'b111011101110;
20'b00101101110011011111: color_data = 12'b111011101110;
20'b00101101110011100000: color_data = 12'b111011101110;
20'b00101101110011100001: color_data = 12'b111011101110;
20'b00101101110011101110: color_data = 12'b111011101110;
20'b00101101110011101111: color_data = 12'b111011101110;
20'b00101101110011110000: color_data = 12'b111011101110;
20'b00101101110011110001: color_data = 12'b111011101110;
20'b00101101110011110010: color_data = 12'b111011101110;
20'b00101101110011110011: color_data = 12'b111011101110;
20'b00101101110011110100: color_data = 12'b111011101110;
20'b00101101110011110101: color_data = 12'b111011101110;
20'b00101101110011110110: color_data = 12'b111011101110;
20'b00101101110011110111: color_data = 12'b111011101110;
20'b00101101110011111001: color_data = 12'b111011101110;
20'b00101101110011111010: color_data = 12'b111011101110;
20'b00101101110011111011: color_data = 12'b111011101110;
20'b00101101110011111100: color_data = 12'b111011101110;
20'b00101101110011111101: color_data = 12'b111011101110;
20'b00101101110011111110: color_data = 12'b111011101110;
20'b00101101110011111111: color_data = 12'b111011101110;
20'b00101101110100000000: color_data = 12'b111011101110;
20'b00101101110100000001: color_data = 12'b111011101110;
20'b00101101110100000010: color_data = 12'b111011101110;
20'b00101101110100100101: color_data = 12'b111011101110;
20'b00101101110100100110: color_data = 12'b111011101110;
20'b00101101110100100111: color_data = 12'b111011101110;
20'b00101101110100101000: color_data = 12'b111011101110;
20'b00101101110100101001: color_data = 12'b111011101110;
20'b00101101110100101010: color_data = 12'b111011101110;
20'b00101101110100101011: color_data = 12'b111011101110;
20'b00101101110100101100: color_data = 12'b111011101110;
20'b00101101110100101101: color_data = 12'b111011101110;
20'b00101101110100101110: color_data = 12'b111011101110;
20'b00101101110100110000: color_data = 12'b111011101110;
20'b00101101110100110001: color_data = 12'b111011101110;
20'b00101101110100110010: color_data = 12'b111011101110;
20'b00101101110100110011: color_data = 12'b111011101110;
20'b00101101110100110100: color_data = 12'b111011101110;
20'b00101101110100110101: color_data = 12'b111011101110;
20'b00101101110100110110: color_data = 12'b111011101110;
20'b00101101110100110111: color_data = 12'b111011101110;
20'b00101101110100111000: color_data = 12'b111011101110;
20'b00101101110100111001: color_data = 12'b111011101110;
20'b00101101110101000110: color_data = 12'b111011101110;
20'b00101101110101000111: color_data = 12'b111011101110;
20'b00101101110101001000: color_data = 12'b111011101110;
20'b00101101110101001001: color_data = 12'b111011101110;
20'b00101101110101001010: color_data = 12'b111011101110;
20'b00101101110101001011: color_data = 12'b111011101110;
20'b00101101110101001100: color_data = 12'b111011101110;
20'b00101101110101001101: color_data = 12'b111011101110;
20'b00101101110101001110: color_data = 12'b111011101110;
20'b00101101110101001111: color_data = 12'b111011101110;
20'b00101101110101010001: color_data = 12'b111011101110;
20'b00101101110101010010: color_data = 12'b111011101110;
20'b00101101110101010011: color_data = 12'b111011101110;
20'b00101101110101010100: color_data = 12'b111011101110;
20'b00101101110101010101: color_data = 12'b111011101110;
20'b00101101110101010110: color_data = 12'b111011101110;
20'b00101101110101010111: color_data = 12'b111011101110;
20'b00101101110101011000: color_data = 12'b111011101110;
20'b00101101110101011001: color_data = 12'b111011101110;
20'b00101101110101011010: color_data = 12'b111011101110;
20'b00101101110101111101: color_data = 12'b111011101110;
20'b00101101110101111110: color_data = 12'b111011101110;
20'b00101101110101111111: color_data = 12'b111011101110;
20'b00101101110110000000: color_data = 12'b111011101110;
20'b00101101110110000001: color_data = 12'b111011101110;
20'b00101101110110000010: color_data = 12'b111011101110;
20'b00101101110110000011: color_data = 12'b111011101110;
20'b00101101110110000100: color_data = 12'b111011101110;
20'b00101101110110000101: color_data = 12'b111011101110;
20'b00101101110110000110: color_data = 12'b111011101110;
20'b00101101110110001000: color_data = 12'b111011101110;
20'b00101101110110001001: color_data = 12'b111011101110;
20'b00101101110110001010: color_data = 12'b111011101110;
20'b00101101110110001011: color_data = 12'b111011101110;
20'b00101101110110001100: color_data = 12'b111011101110;
20'b00101101110110001101: color_data = 12'b111011101110;
20'b00101101110110001110: color_data = 12'b111011101110;
20'b00101101110110001111: color_data = 12'b111011101110;
20'b00101101110110010000: color_data = 12'b111011101110;
20'b00101101110110010001: color_data = 12'b111011101110;
20'b00101101110110011110: color_data = 12'b111011101110;
20'b00101101110110011111: color_data = 12'b111011101110;
20'b00101101110110100000: color_data = 12'b111011101110;
20'b00101101110110100001: color_data = 12'b111011101110;
20'b00101101110110100010: color_data = 12'b111011101110;
20'b00101101110110100011: color_data = 12'b111011101110;
20'b00101101110110100100: color_data = 12'b111011101110;
20'b00101101110110100101: color_data = 12'b111011101110;
20'b00101101110110100110: color_data = 12'b111011101110;
20'b00101101110110100111: color_data = 12'b111011101110;
20'b00101101110110101001: color_data = 12'b111011101110;
20'b00101101110110101010: color_data = 12'b111011101110;
20'b00101101110110101011: color_data = 12'b111011101110;
20'b00101101110110101100: color_data = 12'b111011101110;
20'b00101101110110101101: color_data = 12'b111011101110;
20'b00101101110110101110: color_data = 12'b111011101110;
20'b00101101110110101111: color_data = 12'b111011101110;
20'b00101101110110110000: color_data = 12'b111011101110;
20'b00101101110110110001: color_data = 12'b111011101110;
20'b00101101110110110010: color_data = 12'b111011101110;
20'b00101101110110110100: color_data = 12'b111011101110;
20'b00101101110110110101: color_data = 12'b111011101110;
20'b00101101110110110110: color_data = 12'b111011101110;
20'b00101101110110110111: color_data = 12'b111011101110;
20'b00101101110110111000: color_data = 12'b111011101110;
20'b00101101110110111001: color_data = 12'b111011101110;
20'b00101101110110111010: color_data = 12'b111011101110;
20'b00101101110110111011: color_data = 12'b111011101110;
20'b00101101110110111100: color_data = 12'b111011101110;
20'b00101101110110111101: color_data = 12'b111011101110;
20'b00101101110110111111: color_data = 12'b111011101110;
20'b00101101110111000000: color_data = 12'b111011101110;
20'b00101101110111000001: color_data = 12'b111011101110;
20'b00101101110111000010: color_data = 12'b111011101110;
20'b00101101110111000011: color_data = 12'b111011101110;
20'b00101101110111000100: color_data = 12'b111011101110;
20'b00101101110111000101: color_data = 12'b111011101110;
20'b00101101110111000110: color_data = 12'b111011101110;
20'b00101101110111000111: color_data = 12'b111011101110;
20'b00101101110111001000: color_data = 12'b111011101110;
20'b00101101110111001010: color_data = 12'b111011101110;
20'b00101101110111001011: color_data = 12'b111011101110;
20'b00101101110111001100: color_data = 12'b111011101110;
20'b00101101110111001101: color_data = 12'b111011101110;
20'b00101101110111001110: color_data = 12'b111011101110;
20'b00101101110111001111: color_data = 12'b111011101110;
20'b00101101110111010000: color_data = 12'b111011101110;
20'b00101101110111010001: color_data = 12'b111011101110;
20'b00101101110111010010: color_data = 12'b111011101110;
20'b00101101110111010011: color_data = 12'b111011101110;
20'b00101101110111010101: color_data = 12'b111011101110;
20'b00101101110111010110: color_data = 12'b111011101110;
20'b00101101110111010111: color_data = 12'b111011101110;
20'b00101101110111011000: color_data = 12'b111011101110;
20'b00101101110111011001: color_data = 12'b111011101110;
20'b00101101110111011010: color_data = 12'b111011101110;
20'b00101101110111011011: color_data = 12'b111011101110;
20'b00101101110111011100: color_data = 12'b111011101110;
20'b00101101110111011101: color_data = 12'b111011101110;
20'b00101101110111011110: color_data = 12'b111011101110;
20'b00101101110111100000: color_data = 12'b111011101110;
20'b00101101110111100001: color_data = 12'b111011101110;
20'b00101101110111100010: color_data = 12'b111011101110;
20'b00101101110111100011: color_data = 12'b111011101110;
20'b00101101110111100100: color_data = 12'b111011101110;
20'b00101101110111100101: color_data = 12'b111011101110;
20'b00101101110111100110: color_data = 12'b111011101110;
20'b00101101110111100111: color_data = 12'b111011101110;
20'b00101101110111101000: color_data = 12'b111011101110;
20'b00101101110111101001: color_data = 12'b111011101110;
20'b00101110000010010110: color_data = 12'b111011101110;
20'b00101110000010010111: color_data = 12'b111011101110;
20'b00101110000010011000: color_data = 12'b111011101110;
20'b00101110000010011001: color_data = 12'b111011101110;
20'b00101110000010011010: color_data = 12'b111011101110;
20'b00101110000010011011: color_data = 12'b111011101110;
20'b00101110000010011100: color_data = 12'b111011101110;
20'b00101110000010011101: color_data = 12'b111011101110;
20'b00101110000010011110: color_data = 12'b111011101110;
20'b00101110000010011111: color_data = 12'b111011101110;
20'b00101110000010100001: color_data = 12'b111011101110;
20'b00101110000010100010: color_data = 12'b111011101110;
20'b00101110000010100011: color_data = 12'b111011101110;
20'b00101110000010100100: color_data = 12'b111011101110;
20'b00101110000010100101: color_data = 12'b111011101110;
20'b00101110000010100110: color_data = 12'b111011101110;
20'b00101110000010100111: color_data = 12'b111011101110;
20'b00101110000010101000: color_data = 12'b111011101110;
20'b00101110000010101001: color_data = 12'b111011101110;
20'b00101110000010101010: color_data = 12'b111011101110;
20'b00101110000010101100: color_data = 12'b111011101110;
20'b00101110000010101101: color_data = 12'b111011101110;
20'b00101110000010101110: color_data = 12'b111011101110;
20'b00101110000010101111: color_data = 12'b111011101110;
20'b00101110000010110000: color_data = 12'b111011101110;
20'b00101110000010110001: color_data = 12'b111011101110;
20'b00101110000010110010: color_data = 12'b111011101110;
20'b00101110000010110011: color_data = 12'b111011101110;
20'b00101110000010110100: color_data = 12'b111011101110;
20'b00101110000010110101: color_data = 12'b111011101110;
20'b00101110000010110111: color_data = 12'b111011101110;
20'b00101110000010111000: color_data = 12'b111011101110;
20'b00101110000010111001: color_data = 12'b111011101110;
20'b00101110000010111010: color_data = 12'b111011101110;
20'b00101110000010111011: color_data = 12'b111011101110;
20'b00101110000010111100: color_data = 12'b111011101110;
20'b00101110000010111101: color_data = 12'b111011101110;
20'b00101110000010111110: color_data = 12'b111011101110;
20'b00101110000010111111: color_data = 12'b111011101110;
20'b00101110000011000000: color_data = 12'b111011101110;
20'b00101110000011000010: color_data = 12'b111011101110;
20'b00101110000011000011: color_data = 12'b111011101110;
20'b00101110000011000100: color_data = 12'b111011101110;
20'b00101110000011000101: color_data = 12'b111011101110;
20'b00101110000011000110: color_data = 12'b111011101110;
20'b00101110000011000111: color_data = 12'b111011101110;
20'b00101110000011001000: color_data = 12'b111011101110;
20'b00101110000011001001: color_data = 12'b111011101110;
20'b00101110000011001010: color_data = 12'b111011101110;
20'b00101110000011001011: color_data = 12'b111011101110;
20'b00101110000011001101: color_data = 12'b111011101110;
20'b00101110000011001110: color_data = 12'b111011101110;
20'b00101110000011001111: color_data = 12'b111011101110;
20'b00101110000011010000: color_data = 12'b111011101110;
20'b00101110000011010001: color_data = 12'b111011101110;
20'b00101110000011010010: color_data = 12'b111011101110;
20'b00101110000011010011: color_data = 12'b111011101110;
20'b00101110000011010100: color_data = 12'b111011101110;
20'b00101110000011010101: color_data = 12'b111011101110;
20'b00101110000011010110: color_data = 12'b111011101110;
20'b00101110000011011000: color_data = 12'b111011101110;
20'b00101110000011011001: color_data = 12'b111011101110;
20'b00101110000011011010: color_data = 12'b111011101110;
20'b00101110000011011011: color_data = 12'b111011101110;
20'b00101110000011011100: color_data = 12'b111011101110;
20'b00101110000011011101: color_data = 12'b111011101110;
20'b00101110000011011110: color_data = 12'b111011101110;
20'b00101110000011011111: color_data = 12'b111011101110;
20'b00101110000011100000: color_data = 12'b111011101110;
20'b00101110000011100001: color_data = 12'b111011101110;
20'b00101110000011101110: color_data = 12'b111011101110;
20'b00101110000011101111: color_data = 12'b111011101110;
20'b00101110000011110000: color_data = 12'b111011101110;
20'b00101110000011110001: color_data = 12'b111011101110;
20'b00101110000011110010: color_data = 12'b111011101110;
20'b00101110000011110011: color_data = 12'b111011101110;
20'b00101110000011110100: color_data = 12'b111011101110;
20'b00101110000011110101: color_data = 12'b111011101110;
20'b00101110000011110110: color_data = 12'b111011101110;
20'b00101110000011110111: color_data = 12'b111011101110;
20'b00101110000011111001: color_data = 12'b111011101110;
20'b00101110000011111010: color_data = 12'b111011101110;
20'b00101110000011111011: color_data = 12'b111011101110;
20'b00101110000011111100: color_data = 12'b111011101110;
20'b00101110000011111101: color_data = 12'b111011101110;
20'b00101110000011111110: color_data = 12'b111011101110;
20'b00101110000011111111: color_data = 12'b111011101110;
20'b00101110000100000000: color_data = 12'b111011101110;
20'b00101110000100000001: color_data = 12'b111011101110;
20'b00101110000100000010: color_data = 12'b111011101110;
20'b00101110000100100101: color_data = 12'b111011101110;
20'b00101110000100100110: color_data = 12'b111011101110;
20'b00101110000100100111: color_data = 12'b111011101110;
20'b00101110000100101000: color_data = 12'b111011101110;
20'b00101110000100101001: color_data = 12'b111011101110;
20'b00101110000100101010: color_data = 12'b111011101110;
20'b00101110000100101011: color_data = 12'b111011101110;
20'b00101110000100101100: color_data = 12'b111011101110;
20'b00101110000100101101: color_data = 12'b111011101110;
20'b00101110000100101110: color_data = 12'b111011101110;
20'b00101110000100110000: color_data = 12'b111011101110;
20'b00101110000100110001: color_data = 12'b111011101110;
20'b00101110000100110010: color_data = 12'b111011101110;
20'b00101110000100110011: color_data = 12'b111011101110;
20'b00101110000100110100: color_data = 12'b111011101110;
20'b00101110000100110101: color_data = 12'b111011101110;
20'b00101110000100110110: color_data = 12'b111011101110;
20'b00101110000100110111: color_data = 12'b111011101110;
20'b00101110000100111000: color_data = 12'b111011101110;
20'b00101110000100111001: color_data = 12'b111011101110;
20'b00101110000101000110: color_data = 12'b111011101110;
20'b00101110000101000111: color_data = 12'b111011101110;
20'b00101110000101001000: color_data = 12'b111011101110;
20'b00101110000101001001: color_data = 12'b111011101110;
20'b00101110000101001010: color_data = 12'b111011101110;
20'b00101110000101001011: color_data = 12'b111011101110;
20'b00101110000101001100: color_data = 12'b111011101110;
20'b00101110000101001101: color_data = 12'b111011101110;
20'b00101110000101001110: color_data = 12'b111011101110;
20'b00101110000101001111: color_data = 12'b111011101110;
20'b00101110000101010001: color_data = 12'b111011101110;
20'b00101110000101010010: color_data = 12'b111011101110;
20'b00101110000101010011: color_data = 12'b111011101110;
20'b00101110000101010100: color_data = 12'b111011101110;
20'b00101110000101010101: color_data = 12'b111011101110;
20'b00101110000101010110: color_data = 12'b111011101110;
20'b00101110000101010111: color_data = 12'b111011101110;
20'b00101110000101011000: color_data = 12'b111011101110;
20'b00101110000101011001: color_data = 12'b111011101110;
20'b00101110000101011010: color_data = 12'b111011101110;
20'b00101110000101111101: color_data = 12'b111011101110;
20'b00101110000101111110: color_data = 12'b111011101110;
20'b00101110000101111111: color_data = 12'b111011101110;
20'b00101110000110000000: color_data = 12'b111011101110;
20'b00101110000110000001: color_data = 12'b111011101110;
20'b00101110000110000010: color_data = 12'b111011101110;
20'b00101110000110000011: color_data = 12'b111011101110;
20'b00101110000110000100: color_data = 12'b111011101110;
20'b00101110000110000101: color_data = 12'b111011101110;
20'b00101110000110000110: color_data = 12'b111011101110;
20'b00101110000110001000: color_data = 12'b111011101110;
20'b00101110000110001001: color_data = 12'b111011101110;
20'b00101110000110001010: color_data = 12'b111011101110;
20'b00101110000110001011: color_data = 12'b111011101110;
20'b00101110000110001100: color_data = 12'b111011101110;
20'b00101110000110001101: color_data = 12'b111011101110;
20'b00101110000110001110: color_data = 12'b111011101110;
20'b00101110000110001111: color_data = 12'b111011101110;
20'b00101110000110010000: color_data = 12'b111011101110;
20'b00101110000110010001: color_data = 12'b111011101110;
20'b00101110000110011110: color_data = 12'b111011101110;
20'b00101110000110011111: color_data = 12'b111011101110;
20'b00101110000110100000: color_data = 12'b111011101110;
20'b00101110000110100001: color_data = 12'b111011101110;
20'b00101110000110100010: color_data = 12'b111011101110;
20'b00101110000110100011: color_data = 12'b111011101110;
20'b00101110000110100100: color_data = 12'b111011101110;
20'b00101110000110100101: color_data = 12'b111011101110;
20'b00101110000110100110: color_data = 12'b111011101110;
20'b00101110000110100111: color_data = 12'b111011101110;
20'b00101110000110101001: color_data = 12'b111011101110;
20'b00101110000110101010: color_data = 12'b111011101110;
20'b00101110000110101011: color_data = 12'b111011101110;
20'b00101110000110101100: color_data = 12'b111011101110;
20'b00101110000110101101: color_data = 12'b111011101110;
20'b00101110000110101110: color_data = 12'b111011101110;
20'b00101110000110101111: color_data = 12'b111011101110;
20'b00101110000110110000: color_data = 12'b111011101110;
20'b00101110000110110001: color_data = 12'b111011101110;
20'b00101110000110110010: color_data = 12'b111011101110;
20'b00101110000110110100: color_data = 12'b111011101110;
20'b00101110000110110101: color_data = 12'b111011101110;
20'b00101110000110110110: color_data = 12'b111011101110;
20'b00101110000110110111: color_data = 12'b111011101110;
20'b00101110000110111000: color_data = 12'b111011101110;
20'b00101110000110111001: color_data = 12'b111011101110;
20'b00101110000110111010: color_data = 12'b111011101110;
20'b00101110000110111011: color_data = 12'b111011101110;
20'b00101110000110111100: color_data = 12'b111011101110;
20'b00101110000110111101: color_data = 12'b111011101110;
20'b00101110000110111111: color_data = 12'b111011101110;
20'b00101110000111000000: color_data = 12'b111011101110;
20'b00101110000111000001: color_data = 12'b111011101110;
20'b00101110000111000010: color_data = 12'b111011101110;
20'b00101110000111000011: color_data = 12'b111011101110;
20'b00101110000111000100: color_data = 12'b111011101110;
20'b00101110000111000101: color_data = 12'b111011101110;
20'b00101110000111000110: color_data = 12'b111011101110;
20'b00101110000111000111: color_data = 12'b111011101110;
20'b00101110000111001000: color_data = 12'b111011101110;
20'b00101110000111001010: color_data = 12'b111011101110;
20'b00101110000111001011: color_data = 12'b111011101110;
20'b00101110000111001100: color_data = 12'b111011101110;
20'b00101110000111001101: color_data = 12'b111011101110;
20'b00101110000111001110: color_data = 12'b111011101110;
20'b00101110000111001111: color_data = 12'b111011101110;
20'b00101110000111010000: color_data = 12'b111011101110;
20'b00101110000111010001: color_data = 12'b111011101110;
20'b00101110000111010010: color_data = 12'b111011101110;
20'b00101110000111010011: color_data = 12'b111011101110;
20'b00101110000111010101: color_data = 12'b111011101110;
20'b00101110000111010110: color_data = 12'b111011101110;
20'b00101110000111010111: color_data = 12'b111011101110;
20'b00101110000111011000: color_data = 12'b111011101110;
20'b00101110000111011001: color_data = 12'b111011101110;
20'b00101110000111011010: color_data = 12'b111011101110;
20'b00101110000111011011: color_data = 12'b111011101110;
20'b00101110000111011100: color_data = 12'b111011101110;
20'b00101110000111011101: color_data = 12'b111011101110;
20'b00101110000111011110: color_data = 12'b111011101110;
20'b00101110000111100000: color_data = 12'b111011101110;
20'b00101110000111100001: color_data = 12'b111011101110;
20'b00101110000111100010: color_data = 12'b111011101110;
20'b00101110000111100011: color_data = 12'b111011101110;
20'b00101110000111100100: color_data = 12'b111011101110;
20'b00101110000111100101: color_data = 12'b111011101110;
20'b00101110000111100110: color_data = 12'b111011101110;
20'b00101110000111100111: color_data = 12'b111011101110;
20'b00101110000111101000: color_data = 12'b111011101110;
20'b00101110000111101001: color_data = 12'b111011101110;
20'b00101110010010010110: color_data = 12'b111011101110;
20'b00101110010010010111: color_data = 12'b111011101110;
20'b00101110010010011000: color_data = 12'b111011101110;
20'b00101110010010011001: color_data = 12'b111011101110;
20'b00101110010010011010: color_data = 12'b111011101110;
20'b00101110010010011011: color_data = 12'b111011101110;
20'b00101110010010011100: color_data = 12'b111011101110;
20'b00101110010010011101: color_data = 12'b111011101110;
20'b00101110010010011110: color_data = 12'b111011101110;
20'b00101110010010011111: color_data = 12'b111011101110;
20'b00101110010010100001: color_data = 12'b111011101110;
20'b00101110010010100010: color_data = 12'b111011101110;
20'b00101110010010100011: color_data = 12'b111011101110;
20'b00101110010010100100: color_data = 12'b111011101110;
20'b00101110010010100101: color_data = 12'b111011101110;
20'b00101110010010100110: color_data = 12'b111011101110;
20'b00101110010010100111: color_data = 12'b111011101110;
20'b00101110010010101000: color_data = 12'b111011101110;
20'b00101110010010101001: color_data = 12'b111011101110;
20'b00101110010010101010: color_data = 12'b111011101110;
20'b00101110010010101100: color_data = 12'b111011101110;
20'b00101110010010101101: color_data = 12'b111011101110;
20'b00101110010010101110: color_data = 12'b111011101110;
20'b00101110010010101111: color_data = 12'b111011101110;
20'b00101110010010110000: color_data = 12'b111011101110;
20'b00101110010010110001: color_data = 12'b111011101110;
20'b00101110010010110010: color_data = 12'b111011101110;
20'b00101110010010110011: color_data = 12'b111011101110;
20'b00101110010010110100: color_data = 12'b111011101110;
20'b00101110010010110101: color_data = 12'b111011101110;
20'b00101110010010110111: color_data = 12'b111011101110;
20'b00101110010010111000: color_data = 12'b111011101110;
20'b00101110010010111001: color_data = 12'b111011101110;
20'b00101110010010111010: color_data = 12'b111011101110;
20'b00101110010010111011: color_data = 12'b111011101110;
20'b00101110010010111100: color_data = 12'b111011101110;
20'b00101110010010111101: color_data = 12'b111011101110;
20'b00101110010010111110: color_data = 12'b111011101110;
20'b00101110010010111111: color_data = 12'b111011101110;
20'b00101110010011000000: color_data = 12'b111011101110;
20'b00101110010011000010: color_data = 12'b111011101110;
20'b00101110010011000011: color_data = 12'b111011101110;
20'b00101110010011000100: color_data = 12'b111011101110;
20'b00101110010011000101: color_data = 12'b111011101110;
20'b00101110010011000110: color_data = 12'b111011101110;
20'b00101110010011000111: color_data = 12'b111011101110;
20'b00101110010011001000: color_data = 12'b111011101110;
20'b00101110010011001001: color_data = 12'b111011101110;
20'b00101110010011001010: color_data = 12'b111011101110;
20'b00101110010011001011: color_data = 12'b111011101110;
20'b00101110010011001101: color_data = 12'b111011101110;
20'b00101110010011001110: color_data = 12'b111011101110;
20'b00101110010011001111: color_data = 12'b111011101110;
20'b00101110010011010000: color_data = 12'b111011101110;
20'b00101110010011010001: color_data = 12'b111011101110;
20'b00101110010011010010: color_data = 12'b111011101110;
20'b00101110010011010011: color_data = 12'b111011101110;
20'b00101110010011010100: color_data = 12'b111011101110;
20'b00101110010011010101: color_data = 12'b111011101110;
20'b00101110010011010110: color_data = 12'b111011101110;
20'b00101110010011011000: color_data = 12'b111011101110;
20'b00101110010011011001: color_data = 12'b111011101110;
20'b00101110010011011010: color_data = 12'b111011101110;
20'b00101110010011011011: color_data = 12'b111011101110;
20'b00101110010011011100: color_data = 12'b111011101110;
20'b00101110010011011101: color_data = 12'b111011101110;
20'b00101110010011011110: color_data = 12'b111011101110;
20'b00101110010011011111: color_data = 12'b111011101110;
20'b00101110010011100000: color_data = 12'b111011101110;
20'b00101110010011100001: color_data = 12'b111011101110;
20'b00101110010011101110: color_data = 12'b111011101110;
20'b00101110010011101111: color_data = 12'b111011101110;
20'b00101110010011110000: color_data = 12'b111011101110;
20'b00101110010011110001: color_data = 12'b111011101110;
20'b00101110010011110010: color_data = 12'b111011101110;
20'b00101110010011110011: color_data = 12'b111011101110;
20'b00101110010011110100: color_data = 12'b111011101110;
20'b00101110010011110101: color_data = 12'b111011101110;
20'b00101110010011110110: color_data = 12'b111011101110;
20'b00101110010011110111: color_data = 12'b111011101110;
20'b00101110010011111001: color_data = 12'b111011101110;
20'b00101110010011111010: color_data = 12'b111011101110;
20'b00101110010011111011: color_data = 12'b111011101110;
20'b00101110010011111100: color_data = 12'b111011101110;
20'b00101110010011111101: color_data = 12'b111011101110;
20'b00101110010011111110: color_data = 12'b111011101110;
20'b00101110010011111111: color_data = 12'b111011101110;
20'b00101110010100000000: color_data = 12'b111011101110;
20'b00101110010100000001: color_data = 12'b111011101110;
20'b00101110010100000010: color_data = 12'b111011101110;
20'b00101110010100100101: color_data = 12'b111011101110;
20'b00101110010100100110: color_data = 12'b111011101110;
20'b00101110010100100111: color_data = 12'b111011101110;
20'b00101110010100101000: color_data = 12'b111011101110;
20'b00101110010100101001: color_data = 12'b111011101110;
20'b00101110010100101010: color_data = 12'b111011101110;
20'b00101110010100101011: color_data = 12'b111011101110;
20'b00101110010100101100: color_data = 12'b111011101110;
20'b00101110010100101101: color_data = 12'b111011101110;
20'b00101110010100101110: color_data = 12'b111011101110;
20'b00101110010100110000: color_data = 12'b111011101110;
20'b00101110010100110001: color_data = 12'b111011101110;
20'b00101110010100110010: color_data = 12'b111011101110;
20'b00101110010100110011: color_data = 12'b111011101110;
20'b00101110010100110100: color_data = 12'b111011101110;
20'b00101110010100110101: color_data = 12'b111011101110;
20'b00101110010100110110: color_data = 12'b111011101110;
20'b00101110010100110111: color_data = 12'b111011101110;
20'b00101110010100111000: color_data = 12'b111011101110;
20'b00101110010100111001: color_data = 12'b111011101110;
20'b00101110010101000110: color_data = 12'b111011101110;
20'b00101110010101000111: color_data = 12'b111011101110;
20'b00101110010101001000: color_data = 12'b111011101110;
20'b00101110010101001001: color_data = 12'b111011101110;
20'b00101110010101001010: color_data = 12'b111011101110;
20'b00101110010101001011: color_data = 12'b111011101110;
20'b00101110010101001100: color_data = 12'b111011101110;
20'b00101110010101001101: color_data = 12'b111011101110;
20'b00101110010101001110: color_data = 12'b111011101110;
20'b00101110010101001111: color_data = 12'b111011101110;
20'b00101110010101010001: color_data = 12'b111011101110;
20'b00101110010101010010: color_data = 12'b111011101110;
20'b00101110010101010011: color_data = 12'b111011101110;
20'b00101110010101010100: color_data = 12'b111011101110;
20'b00101110010101010101: color_data = 12'b111011101110;
20'b00101110010101010110: color_data = 12'b111011101110;
20'b00101110010101010111: color_data = 12'b111011101110;
20'b00101110010101011000: color_data = 12'b111011101110;
20'b00101110010101011001: color_data = 12'b111011101110;
20'b00101110010101011010: color_data = 12'b111011101110;
20'b00101110010101111101: color_data = 12'b111011101110;
20'b00101110010101111110: color_data = 12'b111011101110;
20'b00101110010101111111: color_data = 12'b111011101110;
20'b00101110010110000000: color_data = 12'b111011101110;
20'b00101110010110000001: color_data = 12'b111011101110;
20'b00101110010110000010: color_data = 12'b111011101110;
20'b00101110010110000011: color_data = 12'b111011101110;
20'b00101110010110000100: color_data = 12'b111011101110;
20'b00101110010110000101: color_data = 12'b111011101110;
20'b00101110010110000110: color_data = 12'b111011101110;
20'b00101110010110001000: color_data = 12'b111011101110;
20'b00101110010110001001: color_data = 12'b111011101110;
20'b00101110010110001010: color_data = 12'b111011101110;
20'b00101110010110001011: color_data = 12'b111011101110;
20'b00101110010110001100: color_data = 12'b111011101110;
20'b00101110010110001101: color_data = 12'b111011101110;
20'b00101110010110001110: color_data = 12'b111011101110;
20'b00101110010110001111: color_data = 12'b111011101110;
20'b00101110010110010000: color_data = 12'b111011101110;
20'b00101110010110010001: color_data = 12'b111011101110;
20'b00101110010110011110: color_data = 12'b111011101110;
20'b00101110010110011111: color_data = 12'b111011101110;
20'b00101110010110100000: color_data = 12'b111011101110;
20'b00101110010110100001: color_data = 12'b111011101110;
20'b00101110010110100010: color_data = 12'b111011101110;
20'b00101110010110100011: color_data = 12'b111011101110;
20'b00101110010110100100: color_data = 12'b111011101110;
20'b00101110010110100101: color_data = 12'b111011101110;
20'b00101110010110100110: color_data = 12'b111011101110;
20'b00101110010110100111: color_data = 12'b111011101110;
20'b00101110010110101001: color_data = 12'b111011101110;
20'b00101110010110101010: color_data = 12'b111011101110;
20'b00101110010110101011: color_data = 12'b111011101110;
20'b00101110010110101100: color_data = 12'b111011101110;
20'b00101110010110101101: color_data = 12'b111011101110;
20'b00101110010110101110: color_data = 12'b111011101110;
20'b00101110010110101111: color_data = 12'b111011101110;
20'b00101110010110110000: color_data = 12'b111011101110;
20'b00101110010110110001: color_data = 12'b111011101110;
20'b00101110010110110010: color_data = 12'b111011101110;
20'b00101110010110110100: color_data = 12'b111011101110;
20'b00101110010110110101: color_data = 12'b111011101110;
20'b00101110010110110110: color_data = 12'b111011101110;
20'b00101110010110110111: color_data = 12'b111011101110;
20'b00101110010110111000: color_data = 12'b111011101110;
20'b00101110010110111001: color_data = 12'b111011101110;
20'b00101110010110111010: color_data = 12'b111011101110;
20'b00101110010110111011: color_data = 12'b111011101110;
20'b00101110010110111100: color_data = 12'b111011101110;
20'b00101110010110111101: color_data = 12'b111011101110;
20'b00101110010110111111: color_data = 12'b111011101110;
20'b00101110010111000000: color_data = 12'b111011101110;
20'b00101110010111000001: color_data = 12'b111011101110;
20'b00101110010111000010: color_data = 12'b111011101110;
20'b00101110010111000011: color_data = 12'b111011101110;
20'b00101110010111000100: color_data = 12'b111011101110;
20'b00101110010111000101: color_data = 12'b111011101110;
20'b00101110010111000110: color_data = 12'b111011101110;
20'b00101110010111000111: color_data = 12'b111011101110;
20'b00101110010111001000: color_data = 12'b111011101110;
20'b00101110010111001010: color_data = 12'b111011101110;
20'b00101110010111001011: color_data = 12'b111011101110;
20'b00101110010111001100: color_data = 12'b111011101110;
20'b00101110010111001101: color_data = 12'b111011101110;
20'b00101110010111001110: color_data = 12'b111011101110;
20'b00101110010111001111: color_data = 12'b111011101110;
20'b00101110010111010000: color_data = 12'b111011101110;
20'b00101110010111010001: color_data = 12'b111011101110;
20'b00101110010111010010: color_data = 12'b111011101110;
20'b00101110010111010011: color_data = 12'b111011101110;
20'b00101110010111010101: color_data = 12'b111011101110;
20'b00101110010111010110: color_data = 12'b111011101110;
20'b00101110010111010111: color_data = 12'b111011101110;
20'b00101110010111011000: color_data = 12'b111011101110;
20'b00101110010111011001: color_data = 12'b111011101110;
20'b00101110010111011010: color_data = 12'b111011101110;
20'b00101110010111011011: color_data = 12'b111011101110;
20'b00101110010111011100: color_data = 12'b111011101110;
20'b00101110010111011101: color_data = 12'b111011101110;
20'b00101110010111011110: color_data = 12'b111011101110;
20'b00101110010111100000: color_data = 12'b111011101110;
20'b00101110010111100001: color_data = 12'b111011101110;
20'b00101110010111100010: color_data = 12'b111011101110;
20'b00101110010111100011: color_data = 12'b111011101110;
20'b00101110010111100100: color_data = 12'b111011101110;
20'b00101110010111100101: color_data = 12'b111011101110;
20'b00101110010111100110: color_data = 12'b111011101110;
20'b00101110010111100111: color_data = 12'b111011101110;
20'b00101110010111101000: color_data = 12'b111011101110;
20'b00101110010111101001: color_data = 12'b111011101110;
20'b00101110100010010110: color_data = 12'b111011101110;
20'b00101110100010010111: color_data = 12'b111011101110;
20'b00101110100010011000: color_data = 12'b111011101110;
20'b00101110100010011001: color_data = 12'b111011101110;
20'b00101110100010011010: color_data = 12'b111011101110;
20'b00101110100010011011: color_data = 12'b111011101110;
20'b00101110100010011100: color_data = 12'b111011101110;
20'b00101110100010011101: color_data = 12'b111011101110;
20'b00101110100010011110: color_data = 12'b111011101110;
20'b00101110100010011111: color_data = 12'b111011101110;
20'b00101110100010100001: color_data = 12'b111011101110;
20'b00101110100010100010: color_data = 12'b111011101110;
20'b00101110100010100011: color_data = 12'b111011101110;
20'b00101110100010100100: color_data = 12'b111011101110;
20'b00101110100010100101: color_data = 12'b111011101110;
20'b00101110100010100110: color_data = 12'b111011101110;
20'b00101110100010100111: color_data = 12'b111011101110;
20'b00101110100010101000: color_data = 12'b111011101110;
20'b00101110100010101001: color_data = 12'b111011101110;
20'b00101110100010101010: color_data = 12'b111011101110;
20'b00101110100010101100: color_data = 12'b111011101110;
20'b00101110100010101101: color_data = 12'b111011101110;
20'b00101110100010101110: color_data = 12'b111011101110;
20'b00101110100010101111: color_data = 12'b111011101110;
20'b00101110100010110000: color_data = 12'b111011101110;
20'b00101110100010110001: color_data = 12'b111011101110;
20'b00101110100010110010: color_data = 12'b111011101110;
20'b00101110100010110011: color_data = 12'b111011101110;
20'b00101110100010110100: color_data = 12'b111011101110;
20'b00101110100010110101: color_data = 12'b111011101110;
20'b00101110100010110111: color_data = 12'b111011101110;
20'b00101110100010111000: color_data = 12'b111011101110;
20'b00101110100010111001: color_data = 12'b111011101110;
20'b00101110100010111010: color_data = 12'b111011101110;
20'b00101110100010111011: color_data = 12'b111011101110;
20'b00101110100010111100: color_data = 12'b111011101110;
20'b00101110100010111101: color_data = 12'b111011101110;
20'b00101110100010111110: color_data = 12'b111011101110;
20'b00101110100010111111: color_data = 12'b111011101110;
20'b00101110100011000000: color_data = 12'b111011101110;
20'b00101110100011000010: color_data = 12'b111011101110;
20'b00101110100011000011: color_data = 12'b111011101110;
20'b00101110100011000100: color_data = 12'b111011101110;
20'b00101110100011000101: color_data = 12'b111011101110;
20'b00101110100011000110: color_data = 12'b111011101110;
20'b00101110100011000111: color_data = 12'b111011101110;
20'b00101110100011001000: color_data = 12'b111011101110;
20'b00101110100011001001: color_data = 12'b111011101110;
20'b00101110100011001010: color_data = 12'b111011101110;
20'b00101110100011001011: color_data = 12'b111011101110;
20'b00101110100011001101: color_data = 12'b111011101110;
20'b00101110100011001110: color_data = 12'b111011101110;
20'b00101110100011001111: color_data = 12'b111011101110;
20'b00101110100011010000: color_data = 12'b111011101110;
20'b00101110100011010001: color_data = 12'b111011101110;
20'b00101110100011010010: color_data = 12'b111011101110;
20'b00101110100011010011: color_data = 12'b111011101110;
20'b00101110100011010100: color_data = 12'b111011101110;
20'b00101110100011010101: color_data = 12'b111011101110;
20'b00101110100011010110: color_data = 12'b111011101110;
20'b00101110100011011000: color_data = 12'b111011101110;
20'b00101110100011011001: color_data = 12'b111011101110;
20'b00101110100011011010: color_data = 12'b111011101110;
20'b00101110100011011011: color_data = 12'b111011101110;
20'b00101110100011011100: color_data = 12'b111011101110;
20'b00101110100011011101: color_data = 12'b111011101110;
20'b00101110100011011110: color_data = 12'b111011101110;
20'b00101110100011011111: color_data = 12'b111011101110;
20'b00101110100011100000: color_data = 12'b111011101110;
20'b00101110100011100001: color_data = 12'b111011101110;
20'b00101110100011101110: color_data = 12'b111011101110;
20'b00101110100011101111: color_data = 12'b111011101110;
20'b00101110100011110000: color_data = 12'b111011101110;
20'b00101110100011110001: color_data = 12'b111011101110;
20'b00101110100011110010: color_data = 12'b111011101110;
20'b00101110100011110011: color_data = 12'b111011101110;
20'b00101110100011110100: color_data = 12'b111011101110;
20'b00101110100011110101: color_data = 12'b111011101110;
20'b00101110100011110110: color_data = 12'b111011101110;
20'b00101110100011110111: color_data = 12'b111011101110;
20'b00101110100011111001: color_data = 12'b111011101110;
20'b00101110100011111010: color_data = 12'b111011101110;
20'b00101110100011111011: color_data = 12'b111011101110;
20'b00101110100011111100: color_data = 12'b111011101110;
20'b00101110100011111101: color_data = 12'b111011101110;
20'b00101110100011111110: color_data = 12'b111011101110;
20'b00101110100011111111: color_data = 12'b111011101110;
20'b00101110100100000000: color_data = 12'b111011101110;
20'b00101110100100000001: color_data = 12'b111011101110;
20'b00101110100100000010: color_data = 12'b111011101110;
20'b00101110100100100101: color_data = 12'b111011101110;
20'b00101110100100100110: color_data = 12'b111011101110;
20'b00101110100100100111: color_data = 12'b111011101110;
20'b00101110100100101000: color_data = 12'b111011101110;
20'b00101110100100101001: color_data = 12'b111011101110;
20'b00101110100100101010: color_data = 12'b111011101110;
20'b00101110100100101011: color_data = 12'b111011101110;
20'b00101110100100101100: color_data = 12'b111011101110;
20'b00101110100100101101: color_data = 12'b111011101110;
20'b00101110100100101110: color_data = 12'b111011101110;
20'b00101110100100110000: color_data = 12'b111011101110;
20'b00101110100100110001: color_data = 12'b111011101110;
20'b00101110100100110010: color_data = 12'b111011101110;
20'b00101110100100110011: color_data = 12'b111011101110;
20'b00101110100100110100: color_data = 12'b111011101110;
20'b00101110100100110101: color_data = 12'b111011101110;
20'b00101110100100110110: color_data = 12'b111011101110;
20'b00101110100100110111: color_data = 12'b111011101110;
20'b00101110100100111000: color_data = 12'b111011101110;
20'b00101110100100111001: color_data = 12'b111011101110;
20'b00101110100101000110: color_data = 12'b111011101110;
20'b00101110100101000111: color_data = 12'b111011101110;
20'b00101110100101001000: color_data = 12'b111011101110;
20'b00101110100101001001: color_data = 12'b111011101110;
20'b00101110100101001010: color_data = 12'b111011101110;
20'b00101110100101001011: color_data = 12'b111011101110;
20'b00101110100101001100: color_data = 12'b111011101110;
20'b00101110100101001101: color_data = 12'b111011101110;
20'b00101110100101001110: color_data = 12'b111011101110;
20'b00101110100101001111: color_data = 12'b111011101110;
20'b00101110100101010001: color_data = 12'b111011101110;
20'b00101110100101010010: color_data = 12'b111011101110;
20'b00101110100101010011: color_data = 12'b111011101110;
20'b00101110100101010100: color_data = 12'b111011101110;
20'b00101110100101010101: color_data = 12'b111011101110;
20'b00101110100101010110: color_data = 12'b111011101110;
20'b00101110100101010111: color_data = 12'b111011101110;
20'b00101110100101011000: color_data = 12'b111011101110;
20'b00101110100101011001: color_data = 12'b111011101110;
20'b00101110100101011010: color_data = 12'b111011101110;
20'b00101110100101111101: color_data = 12'b111011101110;
20'b00101110100101111110: color_data = 12'b111011101110;
20'b00101110100101111111: color_data = 12'b111011101110;
20'b00101110100110000000: color_data = 12'b111011101110;
20'b00101110100110000001: color_data = 12'b111011101110;
20'b00101110100110000010: color_data = 12'b111011101110;
20'b00101110100110000011: color_data = 12'b111011101110;
20'b00101110100110000100: color_data = 12'b111011101110;
20'b00101110100110000101: color_data = 12'b111011101110;
20'b00101110100110000110: color_data = 12'b111011101110;
20'b00101110100110001000: color_data = 12'b111011101110;
20'b00101110100110001001: color_data = 12'b111011101110;
20'b00101110100110001010: color_data = 12'b111011101110;
20'b00101110100110001011: color_data = 12'b111011101110;
20'b00101110100110001100: color_data = 12'b111011101110;
20'b00101110100110001101: color_data = 12'b111011101110;
20'b00101110100110001110: color_data = 12'b111011101110;
20'b00101110100110001111: color_data = 12'b111011101110;
20'b00101110100110010000: color_data = 12'b111011101110;
20'b00101110100110010001: color_data = 12'b111011101110;
20'b00101110100110011110: color_data = 12'b111011101110;
20'b00101110100110011111: color_data = 12'b111011101110;
20'b00101110100110100000: color_data = 12'b111011101110;
20'b00101110100110100001: color_data = 12'b111011101110;
20'b00101110100110100010: color_data = 12'b111011101110;
20'b00101110100110100011: color_data = 12'b111011101110;
20'b00101110100110100100: color_data = 12'b111011101110;
20'b00101110100110100101: color_data = 12'b111011101110;
20'b00101110100110100110: color_data = 12'b111011101110;
20'b00101110100110100111: color_data = 12'b111011101110;
20'b00101110100110101001: color_data = 12'b111011101110;
20'b00101110100110101010: color_data = 12'b111011101110;
20'b00101110100110101011: color_data = 12'b111011101110;
20'b00101110100110101100: color_data = 12'b111011101110;
20'b00101110100110101101: color_data = 12'b111011101110;
20'b00101110100110101110: color_data = 12'b111011101110;
20'b00101110100110101111: color_data = 12'b111011101110;
20'b00101110100110110000: color_data = 12'b111011101110;
20'b00101110100110110001: color_data = 12'b111011101110;
20'b00101110100110110010: color_data = 12'b111011101110;
20'b00101110100110110100: color_data = 12'b111011101110;
20'b00101110100110110101: color_data = 12'b111011101110;
20'b00101110100110110110: color_data = 12'b111011101110;
20'b00101110100110110111: color_data = 12'b111011101110;
20'b00101110100110111000: color_data = 12'b111011101110;
20'b00101110100110111001: color_data = 12'b111011101110;
20'b00101110100110111010: color_data = 12'b111011101110;
20'b00101110100110111011: color_data = 12'b111011101110;
20'b00101110100110111100: color_data = 12'b111011101110;
20'b00101110100110111101: color_data = 12'b111011101110;
20'b00101110100110111111: color_data = 12'b111011101110;
20'b00101110100111000000: color_data = 12'b111011101110;
20'b00101110100111000001: color_data = 12'b111011101110;
20'b00101110100111000010: color_data = 12'b111011101110;
20'b00101110100111000011: color_data = 12'b111011101110;
20'b00101110100111000100: color_data = 12'b111011101110;
20'b00101110100111000101: color_data = 12'b111011101110;
20'b00101110100111000110: color_data = 12'b111011101110;
20'b00101110100111000111: color_data = 12'b111011101110;
20'b00101110100111001000: color_data = 12'b111011101110;
20'b00101110100111001010: color_data = 12'b111011101110;
20'b00101110100111001011: color_data = 12'b111011101110;
20'b00101110100111001100: color_data = 12'b111011101110;
20'b00101110100111001101: color_data = 12'b111011101110;
20'b00101110100111001110: color_data = 12'b111011101110;
20'b00101110100111001111: color_data = 12'b111011101110;
20'b00101110100111010000: color_data = 12'b111011101110;
20'b00101110100111010001: color_data = 12'b111011101110;
20'b00101110100111010010: color_data = 12'b111011101110;
20'b00101110100111010011: color_data = 12'b111011101110;
20'b00101110100111010101: color_data = 12'b111011101110;
20'b00101110100111010110: color_data = 12'b111011101110;
20'b00101110100111010111: color_data = 12'b111011101110;
20'b00101110100111011000: color_data = 12'b111011101110;
20'b00101110100111011001: color_data = 12'b111011101110;
20'b00101110100111011010: color_data = 12'b111011101110;
20'b00101110100111011011: color_data = 12'b111011101110;
20'b00101110100111011100: color_data = 12'b111011101110;
20'b00101110100111011101: color_data = 12'b111011101110;
20'b00101110100111011110: color_data = 12'b111011101110;
20'b00101110100111100000: color_data = 12'b111011101110;
20'b00101110100111100001: color_data = 12'b111011101110;
20'b00101110100111100010: color_data = 12'b111011101110;
20'b00101110100111100011: color_data = 12'b111011101110;
20'b00101110100111100100: color_data = 12'b111011101110;
20'b00101110100111100101: color_data = 12'b111011101110;
20'b00101110100111100110: color_data = 12'b111011101110;
20'b00101110100111100111: color_data = 12'b111011101110;
20'b00101110100111101000: color_data = 12'b111011101110;
20'b00101110100111101001: color_data = 12'b111011101110;
20'b00101111000010100001: color_data = 12'b111011101110;
20'b00101111000010100010: color_data = 12'b111011101110;
20'b00101111000010100011: color_data = 12'b111011101110;
20'b00101111000010100100: color_data = 12'b111011101110;
20'b00101111000010100101: color_data = 12'b111011101110;
20'b00101111000010100110: color_data = 12'b111011101110;
20'b00101111000010100111: color_data = 12'b111011101110;
20'b00101111000010101000: color_data = 12'b111011101110;
20'b00101111000010101001: color_data = 12'b111011101110;
20'b00101111000010101010: color_data = 12'b111011101110;
20'b00101111000010101100: color_data = 12'b111011101110;
20'b00101111000010101101: color_data = 12'b111011101110;
20'b00101111000010101110: color_data = 12'b111011101110;
20'b00101111000010101111: color_data = 12'b111011101110;
20'b00101111000010110000: color_data = 12'b111011101110;
20'b00101111000010110001: color_data = 12'b111011101110;
20'b00101111000010110010: color_data = 12'b111011101110;
20'b00101111000010110011: color_data = 12'b111011101110;
20'b00101111000010110100: color_data = 12'b111011101110;
20'b00101111000010110101: color_data = 12'b111011101110;
20'b00101111000010110111: color_data = 12'b111011101110;
20'b00101111000010111000: color_data = 12'b111011101110;
20'b00101111000010111001: color_data = 12'b111011101110;
20'b00101111000010111010: color_data = 12'b111011101110;
20'b00101111000010111011: color_data = 12'b111011101110;
20'b00101111000010111100: color_data = 12'b111011101110;
20'b00101111000010111101: color_data = 12'b111011101110;
20'b00101111000010111110: color_data = 12'b111011101110;
20'b00101111000010111111: color_data = 12'b111011101110;
20'b00101111000011000000: color_data = 12'b111011101110;
20'b00101111000011000010: color_data = 12'b111011101110;
20'b00101111000011000011: color_data = 12'b111011101110;
20'b00101111000011000100: color_data = 12'b111011101110;
20'b00101111000011000101: color_data = 12'b111011101110;
20'b00101111000011000110: color_data = 12'b111011101110;
20'b00101111000011000111: color_data = 12'b111011101110;
20'b00101111000011001000: color_data = 12'b111011101110;
20'b00101111000011001001: color_data = 12'b111011101110;
20'b00101111000011001010: color_data = 12'b111011101110;
20'b00101111000011001011: color_data = 12'b111011101110;
20'b00101111000011001101: color_data = 12'b111011101110;
20'b00101111000011001110: color_data = 12'b111011101110;
20'b00101111000011001111: color_data = 12'b111011101110;
20'b00101111000011010000: color_data = 12'b111011101110;
20'b00101111000011010001: color_data = 12'b111011101110;
20'b00101111000011010010: color_data = 12'b111011101110;
20'b00101111000011010011: color_data = 12'b111011101110;
20'b00101111000011010100: color_data = 12'b111011101110;
20'b00101111000011010101: color_data = 12'b111011101110;
20'b00101111000011010110: color_data = 12'b111011101110;
20'b00101111000011101110: color_data = 12'b111011101110;
20'b00101111000011101111: color_data = 12'b111011101110;
20'b00101111000011110000: color_data = 12'b111011101110;
20'b00101111000011110001: color_data = 12'b111011101110;
20'b00101111000011110010: color_data = 12'b111011101110;
20'b00101111000011110011: color_data = 12'b111011101110;
20'b00101111000011110100: color_data = 12'b111011101110;
20'b00101111000011110101: color_data = 12'b111011101110;
20'b00101111000011110110: color_data = 12'b111011101110;
20'b00101111000011110111: color_data = 12'b111011101110;
20'b00101111000011111001: color_data = 12'b111011101110;
20'b00101111000011111010: color_data = 12'b111011101110;
20'b00101111000011111011: color_data = 12'b111011101110;
20'b00101111000011111100: color_data = 12'b111011101110;
20'b00101111000011111101: color_data = 12'b111011101110;
20'b00101111000011111110: color_data = 12'b111011101110;
20'b00101111000011111111: color_data = 12'b111011101110;
20'b00101111000100000000: color_data = 12'b111011101110;
20'b00101111000100000001: color_data = 12'b111011101110;
20'b00101111000100000010: color_data = 12'b111011101110;
20'b00101111000100100101: color_data = 12'b111011101110;
20'b00101111000100100110: color_data = 12'b111011101110;
20'b00101111000100100111: color_data = 12'b111011101110;
20'b00101111000100101000: color_data = 12'b111011101110;
20'b00101111000100101001: color_data = 12'b111011101110;
20'b00101111000100101010: color_data = 12'b111011101110;
20'b00101111000100101011: color_data = 12'b111011101110;
20'b00101111000100101100: color_data = 12'b111011101110;
20'b00101111000100101101: color_data = 12'b111011101110;
20'b00101111000100101110: color_data = 12'b111011101110;
20'b00101111000100110000: color_data = 12'b111011101110;
20'b00101111000100110001: color_data = 12'b111011101110;
20'b00101111000100110010: color_data = 12'b111011101110;
20'b00101111000100110011: color_data = 12'b111011101110;
20'b00101111000100110100: color_data = 12'b111011101110;
20'b00101111000100110101: color_data = 12'b111011101110;
20'b00101111000100110110: color_data = 12'b111011101110;
20'b00101111000100110111: color_data = 12'b111011101110;
20'b00101111000100111000: color_data = 12'b111011101110;
20'b00101111000100111001: color_data = 12'b111011101110;
20'b00101111000101000110: color_data = 12'b111011101110;
20'b00101111000101000111: color_data = 12'b111011101110;
20'b00101111000101001000: color_data = 12'b111011101110;
20'b00101111000101001001: color_data = 12'b111011101110;
20'b00101111000101001010: color_data = 12'b111011101110;
20'b00101111000101001011: color_data = 12'b111011101110;
20'b00101111000101001100: color_data = 12'b111011101110;
20'b00101111000101001101: color_data = 12'b111011101110;
20'b00101111000101001110: color_data = 12'b111011101110;
20'b00101111000101001111: color_data = 12'b111011101110;
20'b00101111000101010001: color_data = 12'b111011101110;
20'b00101111000101010010: color_data = 12'b111011101110;
20'b00101111000101010011: color_data = 12'b111011101110;
20'b00101111000101010100: color_data = 12'b111011101110;
20'b00101111000101010101: color_data = 12'b111011101110;
20'b00101111000101010110: color_data = 12'b111011101110;
20'b00101111000101010111: color_data = 12'b111011101110;
20'b00101111000101011000: color_data = 12'b111011101110;
20'b00101111000101011001: color_data = 12'b111011101110;
20'b00101111000101011010: color_data = 12'b111011101110;
20'b00101111000101111101: color_data = 12'b111011101110;
20'b00101111000101111110: color_data = 12'b111011101110;
20'b00101111000101111111: color_data = 12'b111011101110;
20'b00101111000110000000: color_data = 12'b111011101110;
20'b00101111000110000001: color_data = 12'b111011101110;
20'b00101111000110000010: color_data = 12'b111011101110;
20'b00101111000110000011: color_data = 12'b111011101110;
20'b00101111000110000100: color_data = 12'b111011101110;
20'b00101111000110000101: color_data = 12'b111011101110;
20'b00101111000110000110: color_data = 12'b111011101110;
20'b00101111000110001000: color_data = 12'b111011101110;
20'b00101111000110001001: color_data = 12'b111011101110;
20'b00101111000110001010: color_data = 12'b111011101110;
20'b00101111000110001011: color_data = 12'b111011101110;
20'b00101111000110001100: color_data = 12'b111011101110;
20'b00101111000110001101: color_data = 12'b111011101110;
20'b00101111000110001110: color_data = 12'b111011101110;
20'b00101111000110001111: color_data = 12'b111011101110;
20'b00101111000110010000: color_data = 12'b111011101110;
20'b00101111000110010001: color_data = 12'b111011101110;
20'b00101111000110011110: color_data = 12'b111011101110;
20'b00101111000110011111: color_data = 12'b111011101110;
20'b00101111000110100000: color_data = 12'b111011101110;
20'b00101111000110100001: color_data = 12'b111011101110;
20'b00101111000110100010: color_data = 12'b111011101110;
20'b00101111000110100011: color_data = 12'b111011101110;
20'b00101111000110100100: color_data = 12'b111011101110;
20'b00101111000110100101: color_data = 12'b111011101110;
20'b00101111000110100110: color_data = 12'b111011101110;
20'b00101111000110100111: color_data = 12'b111011101110;
20'b00101111000110101001: color_data = 12'b111011101110;
20'b00101111000110101010: color_data = 12'b111011101110;
20'b00101111000110101011: color_data = 12'b111011101110;
20'b00101111000110101100: color_data = 12'b111011101110;
20'b00101111000110101101: color_data = 12'b111011101110;
20'b00101111000110101110: color_data = 12'b111011101110;
20'b00101111000110101111: color_data = 12'b111011101110;
20'b00101111000110110000: color_data = 12'b111011101110;
20'b00101111000110110001: color_data = 12'b111011101110;
20'b00101111000110110010: color_data = 12'b111011101110;
20'b00101111000110110100: color_data = 12'b111011101110;
20'b00101111000110110101: color_data = 12'b111011101110;
20'b00101111000110110110: color_data = 12'b111011101110;
20'b00101111000110110111: color_data = 12'b111011101110;
20'b00101111000110111000: color_data = 12'b111011101110;
20'b00101111000110111001: color_data = 12'b111011101110;
20'b00101111000110111010: color_data = 12'b111011101110;
20'b00101111000110111011: color_data = 12'b111011101110;
20'b00101111000110111100: color_data = 12'b111011101110;
20'b00101111000110111101: color_data = 12'b111011101110;
20'b00101111000110111111: color_data = 12'b111011101110;
20'b00101111000111000000: color_data = 12'b111011101110;
20'b00101111000111000001: color_data = 12'b111011101110;
20'b00101111000111000010: color_data = 12'b111011101110;
20'b00101111000111000011: color_data = 12'b111011101110;
20'b00101111000111000100: color_data = 12'b111011101110;
20'b00101111000111000101: color_data = 12'b111011101110;
20'b00101111000111000110: color_data = 12'b111011101110;
20'b00101111000111000111: color_data = 12'b111011101110;
20'b00101111000111001000: color_data = 12'b111011101110;
20'b00101111000111001010: color_data = 12'b111011101110;
20'b00101111000111001011: color_data = 12'b111011101110;
20'b00101111000111001100: color_data = 12'b111011101110;
20'b00101111000111001101: color_data = 12'b111011101110;
20'b00101111000111001110: color_data = 12'b111011101110;
20'b00101111000111001111: color_data = 12'b111011101110;
20'b00101111000111010000: color_data = 12'b111011101110;
20'b00101111000111010001: color_data = 12'b111011101110;
20'b00101111000111010010: color_data = 12'b111011101110;
20'b00101111000111010011: color_data = 12'b111011101110;
20'b00101111000111010101: color_data = 12'b111011101110;
20'b00101111000111010110: color_data = 12'b111011101110;
20'b00101111000111010111: color_data = 12'b111011101110;
20'b00101111000111011000: color_data = 12'b111011101110;
20'b00101111000111011001: color_data = 12'b111011101110;
20'b00101111000111011010: color_data = 12'b111011101110;
20'b00101111000111011011: color_data = 12'b111011101110;
20'b00101111000111011100: color_data = 12'b111011101110;
20'b00101111000111011101: color_data = 12'b111011101110;
20'b00101111000111011110: color_data = 12'b111011101110;
20'b00101111000111100000: color_data = 12'b111011101110;
20'b00101111000111100001: color_data = 12'b111011101110;
20'b00101111000111100010: color_data = 12'b111011101110;
20'b00101111000111100011: color_data = 12'b111011101110;
20'b00101111000111100100: color_data = 12'b111011101110;
20'b00101111000111100101: color_data = 12'b111011101110;
20'b00101111000111100110: color_data = 12'b111011101110;
20'b00101111000111100111: color_data = 12'b111011101110;
20'b00101111000111101000: color_data = 12'b111011101110;
20'b00101111000111101001: color_data = 12'b111011101110;
20'b00101111010010100001: color_data = 12'b111011101110;
20'b00101111010010100010: color_data = 12'b111011101110;
20'b00101111010010100011: color_data = 12'b111011101110;
20'b00101111010010100100: color_data = 12'b111011101110;
20'b00101111010010100101: color_data = 12'b111011101110;
20'b00101111010010100110: color_data = 12'b111011101110;
20'b00101111010010100111: color_data = 12'b111011101110;
20'b00101111010010101000: color_data = 12'b111011101110;
20'b00101111010010101001: color_data = 12'b111011101110;
20'b00101111010010101010: color_data = 12'b111011101110;
20'b00101111010010101100: color_data = 12'b111011101110;
20'b00101111010010101101: color_data = 12'b111011101110;
20'b00101111010010101110: color_data = 12'b111011101110;
20'b00101111010010101111: color_data = 12'b111011101110;
20'b00101111010010110000: color_data = 12'b111011101110;
20'b00101111010010110001: color_data = 12'b111011101110;
20'b00101111010010110010: color_data = 12'b111011101110;
20'b00101111010010110011: color_data = 12'b111011101110;
20'b00101111010010110100: color_data = 12'b111011101110;
20'b00101111010010110101: color_data = 12'b111011101110;
20'b00101111010010110111: color_data = 12'b111011101110;
20'b00101111010010111000: color_data = 12'b111011101110;
20'b00101111010010111001: color_data = 12'b111011101110;
20'b00101111010010111010: color_data = 12'b111011101110;
20'b00101111010010111011: color_data = 12'b111011101110;
20'b00101111010010111100: color_data = 12'b111011101110;
20'b00101111010010111101: color_data = 12'b111011101110;
20'b00101111010010111110: color_data = 12'b111011101110;
20'b00101111010010111111: color_data = 12'b111011101110;
20'b00101111010011000000: color_data = 12'b111011101110;
20'b00101111010011000010: color_data = 12'b111011101110;
20'b00101111010011000011: color_data = 12'b111011101110;
20'b00101111010011000100: color_data = 12'b111011101110;
20'b00101111010011000101: color_data = 12'b111011101110;
20'b00101111010011000110: color_data = 12'b111011101110;
20'b00101111010011000111: color_data = 12'b111011101110;
20'b00101111010011001000: color_data = 12'b111011101110;
20'b00101111010011001001: color_data = 12'b111011101110;
20'b00101111010011001010: color_data = 12'b111011101110;
20'b00101111010011001011: color_data = 12'b111011101110;
20'b00101111010011001101: color_data = 12'b111011101110;
20'b00101111010011001110: color_data = 12'b111011101110;
20'b00101111010011001111: color_data = 12'b111011101110;
20'b00101111010011010000: color_data = 12'b111011101110;
20'b00101111010011010001: color_data = 12'b111011101110;
20'b00101111010011010010: color_data = 12'b111011101110;
20'b00101111010011010011: color_data = 12'b111011101110;
20'b00101111010011010100: color_data = 12'b111011101110;
20'b00101111010011010101: color_data = 12'b111011101110;
20'b00101111010011010110: color_data = 12'b111011101110;
20'b00101111010011101110: color_data = 12'b111011101110;
20'b00101111010011101111: color_data = 12'b111011101110;
20'b00101111010011110000: color_data = 12'b111011101110;
20'b00101111010011110001: color_data = 12'b111011101110;
20'b00101111010011110010: color_data = 12'b111011101110;
20'b00101111010011110011: color_data = 12'b111011101110;
20'b00101111010011110100: color_data = 12'b111011101110;
20'b00101111010011110101: color_data = 12'b111011101110;
20'b00101111010011110110: color_data = 12'b111011101110;
20'b00101111010011110111: color_data = 12'b111011101110;
20'b00101111010011111001: color_data = 12'b111011101110;
20'b00101111010011111010: color_data = 12'b111011101110;
20'b00101111010011111011: color_data = 12'b111011101110;
20'b00101111010011111100: color_data = 12'b111011101110;
20'b00101111010011111101: color_data = 12'b111011101110;
20'b00101111010011111110: color_data = 12'b111011101110;
20'b00101111010011111111: color_data = 12'b111011101110;
20'b00101111010100000000: color_data = 12'b111011101110;
20'b00101111010100000001: color_data = 12'b111011101110;
20'b00101111010100000010: color_data = 12'b111011101110;
20'b00101111010100100101: color_data = 12'b111011101110;
20'b00101111010100100110: color_data = 12'b111011101110;
20'b00101111010100100111: color_data = 12'b111011101110;
20'b00101111010100101000: color_data = 12'b111011101110;
20'b00101111010100101001: color_data = 12'b111011101110;
20'b00101111010100101010: color_data = 12'b111011101110;
20'b00101111010100101011: color_data = 12'b111011101110;
20'b00101111010100101100: color_data = 12'b111011101110;
20'b00101111010100101101: color_data = 12'b111011101110;
20'b00101111010100101110: color_data = 12'b111011101110;
20'b00101111010100110000: color_data = 12'b111011101110;
20'b00101111010100110001: color_data = 12'b111011101110;
20'b00101111010100110010: color_data = 12'b111011101110;
20'b00101111010100110011: color_data = 12'b111011101110;
20'b00101111010100110100: color_data = 12'b111011101110;
20'b00101111010100110101: color_data = 12'b111011101110;
20'b00101111010100110110: color_data = 12'b111011101110;
20'b00101111010100110111: color_data = 12'b111011101110;
20'b00101111010100111000: color_data = 12'b111011101110;
20'b00101111010100111001: color_data = 12'b111011101110;
20'b00101111010101000110: color_data = 12'b111011101110;
20'b00101111010101000111: color_data = 12'b111011101110;
20'b00101111010101001000: color_data = 12'b111011101110;
20'b00101111010101001001: color_data = 12'b111011101110;
20'b00101111010101001010: color_data = 12'b111011101110;
20'b00101111010101001011: color_data = 12'b111011101110;
20'b00101111010101001100: color_data = 12'b111011101110;
20'b00101111010101001101: color_data = 12'b111011101110;
20'b00101111010101001110: color_data = 12'b111011101110;
20'b00101111010101001111: color_data = 12'b111011101110;
20'b00101111010101010001: color_data = 12'b111011101110;
20'b00101111010101010010: color_data = 12'b111011101110;
20'b00101111010101010011: color_data = 12'b111011101110;
20'b00101111010101010100: color_data = 12'b111011101110;
20'b00101111010101010101: color_data = 12'b111011101110;
20'b00101111010101010110: color_data = 12'b111011101110;
20'b00101111010101010111: color_data = 12'b111011101110;
20'b00101111010101011000: color_data = 12'b111011101110;
20'b00101111010101011001: color_data = 12'b111011101110;
20'b00101111010101011010: color_data = 12'b111011101110;
20'b00101111010101111101: color_data = 12'b111011101110;
20'b00101111010101111110: color_data = 12'b111011101110;
20'b00101111010101111111: color_data = 12'b111011101110;
20'b00101111010110000000: color_data = 12'b111011101110;
20'b00101111010110000001: color_data = 12'b111011101110;
20'b00101111010110000010: color_data = 12'b111011101110;
20'b00101111010110000011: color_data = 12'b111011101110;
20'b00101111010110000100: color_data = 12'b111011101110;
20'b00101111010110000101: color_data = 12'b111011101110;
20'b00101111010110000110: color_data = 12'b111011101110;
20'b00101111010110001000: color_data = 12'b111011101110;
20'b00101111010110001001: color_data = 12'b111011101110;
20'b00101111010110001010: color_data = 12'b111011101110;
20'b00101111010110001011: color_data = 12'b111011101110;
20'b00101111010110001100: color_data = 12'b111011101110;
20'b00101111010110001101: color_data = 12'b111011101110;
20'b00101111010110001110: color_data = 12'b111011101110;
20'b00101111010110001111: color_data = 12'b111011101110;
20'b00101111010110010000: color_data = 12'b111011101110;
20'b00101111010110010001: color_data = 12'b111011101110;
20'b00101111010110011110: color_data = 12'b111011101110;
20'b00101111010110011111: color_data = 12'b111011101110;
20'b00101111010110100000: color_data = 12'b111011101110;
20'b00101111010110100001: color_data = 12'b111011101110;
20'b00101111010110100010: color_data = 12'b111011101110;
20'b00101111010110100011: color_data = 12'b111011101110;
20'b00101111010110100100: color_data = 12'b111011101110;
20'b00101111010110100101: color_data = 12'b111011101110;
20'b00101111010110100110: color_data = 12'b111011101110;
20'b00101111010110100111: color_data = 12'b111011101110;
20'b00101111010110101001: color_data = 12'b111011101110;
20'b00101111010110101010: color_data = 12'b111011101110;
20'b00101111010110101011: color_data = 12'b111011101110;
20'b00101111010110101100: color_data = 12'b111011101110;
20'b00101111010110101101: color_data = 12'b111011101110;
20'b00101111010110101110: color_data = 12'b111011101110;
20'b00101111010110101111: color_data = 12'b111011101110;
20'b00101111010110110000: color_data = 12'b111011101110;
20'b00101111010110110001: color_data = 12'b111011101110;
20'b00101111010110110010: color_data = 12'b111011101110;
20'b00101111010110110100: color_data = 12'b111011101110;
20'b00101111010110110101: color_data = 12'b111011101110;
20'b00101111010110110110: color_data = 12'b111011101110;
20'b00101111010110110111: color_data = 12'b111011101110;
20'b00101111010110111000: color_data = 12'b111011101110;
20'b00101111010110111001: color_data = 12'b111011101110;
20'b00101111010110111010: color_data = 12'b111011101110;
20'b00101111010110111011: color_data = 12'b111011101110;
20'b00101111010110111100: color_data = 12'b111011101110;
20'b00101111010110111101: color_data = 12'b111011101110;
20'b00101111010110111111: color_data = 12'b111011101110;
20'b00101111010111000000: color_data = 12'b111011101110;
20'b00101111010111000001: color_data = 12'b111011101110;
20'b00101111010111000010: color_data = 12'b111011101110;
20'b00101111010111000011: color_data = 12'b111011101110;
20'b00101111010111000100: color_data = 12'b111011101110;
20'b00101111010111000101: color_data = 12'b111011101110;
20'b00101111010111000110: color_data = 12'b111011101110;
20'b00101111010111000111: color_data = 12'b111011101110;
20'b00101111010111001000: color_data = 12'b111011101110;
20'b00101111010111001010: color_data = 12'b111011101110;
20'b00101111010111001011: color_data = 12'b111011101110;
20'b00101111010111001100: color_data = 12'b111011101110;
20'b00101111010111001101: color_data = 12'b111011101110;
20'b00101111010111001110: color_data = 12'b111011101110;
20'b00101111010111001111: color_data = 12'b111011101110;
20'b00101111010111010000: color_data = 12'b111011101110;
20'b00101111010111010001: color_data = 12'b111011101110;
20'b00101111010111010010: color_data = 12'b111011101110;
20'b00101111010111010011: color_data = 12'b111011101110;
20'b00101111010111010101: color_data = 12'b111011101110;
20'b00101111010111010110: color_data = 12'b111011101110;
20'b00101111010111010111: color_data = 12'b111011101110;
20'b00101111010111011000: color_data = 12'b111011101110;
20'b00101111010111011001: color_data = 12'b111011101110;
20'b00101111010111011010: color_data = 12'b111011101110;
20'b00101111010111011011: color_data = 12'b111011101110;
20'b00101111010111011100: color_data = 12'b111011101110;
20'b00101111010111011101: color_data = 12'b111011101110;
20'b00101111010111011110: color_data = 12'b111011101110;
20'b00101111010111100000: color_data = 12'b111011101110;
20'b00101111010111100001: color_data = 12'b111011101110;
20'b00101111010111100010: color_data = 12'b111011101110;
20'b00101111010111100011: color_data = 12'b111011101110;
20'b00101111010111100100: color_data = 12'b111011101110;
20'b00101111010111100101: color_data = 12'b111011101110;
20'b00101111010111100110: color_data = 12'b111011101110;
20'b00101111010111100111: color_data = 12'b111011101110;
20'b00101111010111101000: color_data = 12'b111011101110;
20'b00101111010111101001: color_data = 12'b111011101110;
20'b00101111100010100001: color_data = 12'b111011101110;
20'b00101111100010100010: color_data = 12'b111011101110;
20'b00101111100010100011: color_data = 12'b111011101110;
20'b00101111100010100100: color_data = 12'b111011101110;
20'b00101111100010100101: color_data = 12'b111011101110;
20'b00101111100010100110: color_data = 12'b111011101110;
20'b00101111100010100111: color_data = 12'b111011101110;
20'b00101111100010101000: color_data = 12'b111011101110;
20'b00101111100010101001: color_data = 12'b111011101110;
20'b00101111100010101010: color_data = 12'b111011101110;
20'b00101111100010101100: color_data = 12'b111011101110;
20'b00101111100010101101: color_data = 12'b111011101110;
20'b00101111100010101110: color_data = 12'b111011101110;
20'b00101111100010101111: color_data = 12'b111011101110;
20'b00101111100010110000: color_data = 12'b111011101110;
20'b00101111100010110001: color_data = 12'b111011101110;
20'b00101111100010110010: color_data = 12'b111011101110;
20'b00101111100010110011: color_data = 12'b111011101110;
20'b00101111100010110100: color_data = 12'b111011101110;
20'b00101111100010110101: color_data = 12'b111011101110;
20'b00101111100010110111: color_data = 12'b111011101110;
20'b00101111100010111000: color_data = 12'b111011101110;
20'b00101111100010111001: color_data = 12'b111011101110;
20'b00101111100010111010: color_data = 12'b111011101110;
20'b00101111100010111011: color_data = 12'b111011101110;
20'b00101111100010111100: color_data = 12'b111011101110;
20'b00101111100010111101: color_data = 12'b111011101110;
20'b00101111100010111110: color_data = 12'b111011101110;
20'b00101111100010111111: color_data = 12'b111011101110;
20'b00101111100011000000: color_data = 12'b111011101110;
20'b00101111100011000010: color_data = 12'b111011101110;
20'b00101111100011000011: color_data = 12'b111011101110;
20'b00101111100011000100: color_data = 12'b111011101110;
20'b00101111100011000101: color_data = 12'b111011101110;
20'b00101111100011000110: color_data = 12'b111011101110;
20'b00101111100011000111: color_data = 12'b111011101110;
20'b00101111100011001000: color_data = 12'b111011101110;
20'b00101111100011001001: color_data = 12'b111011101110;
20'b00101111100011001010: color_data = 12'b111011101110;
20'b00101111100011001011: color_data = 12'b111011101110;
20'b00101111100011001101: color_data = 12'b111011101110;
20'b00101111100011001110: color_data = 12'b111011101110;
20'b00101111100011001111: color_data = 12'b111011101110;
20'b00101111100011010000: color_data = 12'b111011101110;
20'b00101111100011010001: color_data = 12'b111011101110;
20'b00101111100011010010: color_data = 12'b111011101110;
20'b00101111100011010011: color_data = 12'b111011101110;
20'b00101111100011010100: color_data = 12'b111011101110;
20'b00101111100011010101: color_data = 12'b111011101110;
20'b00101111100011010110: color_data = 12'b111011101110;
20'b00101111100011101110: color_data = 12'b111011101110;
20'b00101111100011101111: color_data = 12'b111011101110;
20'b00101111100011110000: color_data = 12'b111011101110;
20'b00101111100011110001: color_data = 12'b111011101110;
20'b00101111100011110010: color_data = 12'b111011101110;
20'b00101111100011110011: color_data = 12'b111011101110;
20'b00101111100011110100: color_data = 12'b111011101110;
20'b00101111100011110101: color_data = 12'b111011101110;
20'b00101111100011110110: color_data = 12'b111011101110;
20'b00101111100011110111: color_data = 12'b111011101110;
20'b00101111100011111001: color_data = 12'b111011101110;
20'b00101111100011111010: color_data = 12'b111011101110;
20'b00101111100011111011: color_data = 12'b111011101110;
20'b00101111100011111100: color_data = 12'b111011101110;
20'b00101111100011111101: color_data = 12'b111011101110;
20'b00101111100011111110: color_data = 12'b111011101110;
20'b00101111100011111111: color_data = 12'b111011101110;
20'b00101111100100000000: color_data = 12'b111011101110;
20'b00101111100100000001: color_data = 12'b111011101110;
20'b00101111100100000010: color_data = 12'b111011101110;
20'b00101111100100100101: color_data = 12'b111011101110;
20'b00101111100100100110: color_data = 12'b111011101110;
20'b00101111100100100111: color_data = 12'b111011101110;
20'b00101111100100101000: color_data = 12'b111011101110;
20'b00101111100100101001: color_data = 12'b111011101110;
20'b00101111100100101010: color_data = 12'b111011101110;
20'b00101111100100101011: color_data = 12'b111011101110;
20'b00101111100100101100: color_data = 12'b111011101110;
20'b00101111100100101101: color_data = 12'b111011101110;
20'b00101111100100101110: color_data = 12'b111011101110;
20'b00101111100100110000: color_data = 12'b111011101110;
20'b00101111100100110001: color_data = 12'b111011101110;
20'b00101111100100110010: color_data = 12'b111011101110;
20'b00101111100100110011: color_data = 12'b111011101110;
20'b00101111100100110100: color_data = 12'b111011101110;
20'b00101111100100110101: color_data = 12'b111011101110;
20'b00101111100100110110: color_data = 12'b111011101110;
20'b00101111100100110111: color_data = 12'b111011101110;
20'b00101111100100111000: color_data = 12'b111011101110;
20'b00101111100100111001: color_data = 12'b111011101110;
20'b00101111100101000110: color_data = 12'b111011101110;
20'b00101111100101000111: color_data = 12'b111011101110;
20'b00101111100101001000: color_data = 12'b111011101110;
20'b00101111100101001001: color_data = 12'b111011101110;
20'b00101111100101001010: color_data = 12'b111011101110;
20'b00101111100101001011: color_data = 12'b111011101110;
20'b00101111100101001100: color_data = 12'b111011101110;
20'b00101111100101001101: color_data = 12'b111011101110;
20'b00101111100101001110: color_data = 12'b111011101110;
20'b00101111100101001111: color_data = 12'b111011101110;
20'b00101111100101010001: color_data = 12'b111011101110;
20'b00101111100101010010: color_data = 12'b111011101110;
20'b00101111100101010011: color_data = 12'b111011101110;
20'b00101111100101010100: color_data = 12'b111011101110;
20'b00101111100101010101: color_data = 12'b111011101110;
20'b00101111100101010110: color_data = 12'b111011101110;
20'b00101111100101010111: color_data = 12'b111011101110;
20'b00101111100101011000: color_data = 12'b111011101110;
20'b00101111100101011001: color_data = 12'b111011101110;
20'b00101111100101011010: color_data = 12'b111011101110;
20'b00101111100101111101: color_data = 12'b111011101110;
20'b00101111100101111110: color_data = 12'b111011101110;
20'b00101111100101111111: color_data = 12'b111011101110;
20'b00101111100110000000: color_data = 12'b111011101110;
20'b00101111100110000001: color_data = 12'b111011101110;
20'b00101111100110000010: color_data = 12'b111011101110;
20'b00101111100110000011: color_data = 12'b111011101110;
20'b00101111100110000100: color_data = 12'b111011101110;
20'b00101111100110000101: color_data = 12'b111011101110;
20'b00101111100110000110: color_data = 12'b111011101110;
20'b00101111100110001000: color_data = 12'b111011101110;
20'b00101111100110001001: color_data = 12'b111011101110;
20'b00101111100110001010: color_data = 12'b111011101110;
20'b00101111100110001011: color_data = 12'b111011101110;
20'b00101111100110001100: color_data = 12'b111011101110;
20'b00101111100110001101: color_data = 12'b111011101110;
20'b00101111100110001110: color_data = 12'b111011101110;
20'b00101111100110001111: color_data = 12'b111011101110;
20'b00101111100110010000: color_data = 12'b111011101110;
20'b00101111100110010001: color_data = 12'b111011101110;
20'b00101111100110011110: color_data = 12'b111011101110;
20'b00101111100110011111: color_data = 12'b111011101110;
20'b00101111100110100000: color_data = 12'b111011101110;
20'b00101111100110100001: color_data = 12'b111011101110;
20'b00101111100110100010: color_data = 12'b111011101110;
20'b00101111100110100011: color_data = 12'b111011101110;
20'b00101111100110100100: color_data = 12'b111011101110;
20'b00101111100110100101: color_data = 12'b111011101110;
20'b00101111100110100110: color_data = 12'b111011101110;
20'b00101111100110100111: color_data = 12'b111011101110;
20'b00101111100110101001: color_data = 12'b111011101110;
20'b00101111100110101010: color_data = 12'b111011101110;
20'b00101111100110101011: color_data = 12'b111011101110;
20'b00101111100110101100: color_data = 12'b111011101110;
20'b00101111100110101101: color_data = 12'b111011101110;
20'b00101111100110101110: color_data = 12'b111011101110;
20'b00101111100110101111: color_data = 12'b111011101110;
20'b00101111100110110000: color_data = 12'b111011101110;
20'b00101111100110110001: color_data = 12'b111011101110;
20'b00101111100110110010: color_data = 12'b111011101110;
20'b00101111100110110100: color_data = 12'b111011101110;
20'b00101111100110110101: color_data = 12'b111011101110;
20'b00101111100110110110: color_data = 12'b111011101110;
20'b00101111100110110111: color_data = 12'b111011101110;
20'b00101111100110111000: color_data = 12'b111011101110;
20'b00101111100110111001: color_data = 12'b111011101110;
20'b00101111100110111010: color_data = 12'b111011101110;
20'b00101111100110111011: color_data = 12'b111011101110;
20'b00101111100110111100: color_data = 12'b111011101110;
20'b00101111100110111101: color_data = 12'b111011101110;
20'b00101111100110111111: color_data = 12'b111011101110;
20'b00101111100111000000: color_data = 12'b111011101110;
20'b00101111100111000001: color_data = 12'b111011101110;
20'b00101111100111000010: color_data = 12'b111011101110;
20'b00101111100111000011: color_data = 12'b111011101110;
20'b00101111100111000100: color_data = 12'b111011101110;
20'b00101111100111000101: color_data = 12'b111011101110;
20'b00101111100111000110: color_data = 12'b111011101110;
20'b00101111100111000111: color_data = 12'b111011101110;
20'b00101111100111001000: color_data = 12'b111011101110;
20'b00101111100111001010: color_data = 12'b111011101110;
20'b00101111100111001011: color_data = 12'b111011101110;
20'b00101111100111001100: color_data = 12'b111011101110;
20'b00101111100111001101: color_data = 12'b111011101110;
20'b00101111100111001110: color_data = 12'b111011101110;
20'b00101111100111001111: color_data = 12'b111011101110;
20'b00101111100111010000: color_data = 12'b111011101110;
20'b00101111100111010001: color_data = 12'b111011101110;
20'b00101111100111010010: color_data = 12'b111011101110;
20'b00101111100111010011: color_data = 12'b111011101110;
20'b00101111100111010101: color_data = 12'b111011101110;
20'b00101111100111010110: color_data = 12'b111011101110;
20'b00101111100111010111: color_data = 12'b111011101110;
20'b00101111100111011000: color_data = 12'b111011101110;
20'b00101111100111011001: color_data = 12'b111011101110;
20'b00101111100111011010: color_data = 12'b111011101110;
20'b00101111100111011011: color_data = 12'b111011101110;
20'b00101111100111011100: color_data = 12'b111011101110;
20'b00101111100111011101: color_data = 12'b111011101110;
20'b00101111100111011110: color_data = 12'b111011101110;
20'b00101111100111100000: color_data = 12'b111011101110;
20'b00101111100111100001: color_data = 12'b111011101110;
20'b00101111100111100010: color_data = 12'b111011101110;
20'b00101111100111100011: color_data = 12'b111011101110;
20'b00101111100111100100: color_data = 12'b111011101110;
20'b00101111100111100101: color_data = 12'b111011101110;
20'b00101111100111100110: color_data = 12'b111011101110;
20'b00101111100111100111: color_data = 12'b111011101110;
20'b00101111100111101000: color_data = 12'b111011101110;
20'b00101111100111101001: color_data = 12'b111011101110;
20'b00101111110010100001: color_data = 12'b111011101110;
20'b00101111110010100010: color_data = 12'b111011101110;
20'b00101111110010100011: color_data = 12'b111011101110;
20'b00101111110010100100: color_data = 12'b111011101110;
20'b00101111110010100101: color_data = 12'b111011101110;
20'b00101111110010100110: color_data = 12'b111011101110;
20'b00101111110010100111: color_data = 12'b111011101110;
20'b00101111110010101000: color_data = 12'b111011101110;
20'b00101111110010101001: color_data = 12'b111011101110;
20'b00101111110010101010: color_data = 12'b111011101110;
20'b00101111110010101100: color_data = 12'b111011101110;
20'b00101111110010101101: color_data = 12'b111011101110;
20'b00101111110010101110: color_data = 12'b111011101110;
20'b00101111110010101111: color_data = 12'b111011101110;
20'b00101111110010110000: color_data = 12'b111011101110;
20'b00101111110010110001: color_data = 12'b111011101110;
20'b00101111110010110010: color_data = 12'b111011101110;
20'b00101111110010110011: color_data = 12'b111011101110;
20'b00101111110010110100: color_data = 12'b111011101110;
20'b00101111110010110101: color_data = 12'b111011101110;
20'b00101111110010110111: color_data = 12'b111011101110;
20'b00101111110010111000: color_data = 12'b111011101110;
20'b00101111110010111001: color_data = 12'b111011101110;
20'b00101111110010111010: color_data = 12'b111011101110;
20'b00101111110010111011: color_data = 12'b111011101110;
20'b00101111110010111100: color_data = 12'b111011101110;
20'b00101111110010111101: color_data = 12'b111011101110;
20'b00101111110010111110: color_data = 12'b111011101110;
20'b00101111110010111111: color_data = 12'b111011101110;
20'b00101111110011000000: color_data = 12'b111011101110;
20'b00101111110011000010: color_data = 12'b111011101110;
20'b00101111110011000011: color_data = 12'b111011101110;
20'b00101111110011000100: color_data = 12'b111011101110;
20'b00101111110011000101: color_data = 12'b111011101110;
20'b00101111110011000110: color_data = 12'b111011101110;
20'b00101111110011000111: color_data = 12'b111011101110;
20'b00101111110011001000: color_data = 12'b111011101110;
20'b00101111110011001001: color_data = 12'b111011101110;
20'b00101111110011001010: color_data = 12'b111011101110;
20'b00101111110011001011: color_data = 12'b111011101110;
20'b00101111110011001101: color_data = 12'b111011101110;
20'b00101111110011001110: color_data = 12'b111011101110;
20'b00101111110011001111: color_data = 12'b111011101110;
20'b00101111110011010000: color_data = 12'b111011101110;
20'b00101111110011010001: color_data = 12'b111011101110;
20'b00101111110011010010: color_data = 12'b111011101110;
20'b00101111110011010011: color_data = 12'b111011101110;
20'b00101111110011010100: color_data = 12'b111011101110;
20'b00101111110011010101: color_data = 12'b111011101110;
20'b00101111110011010110: color_data = 12'b111011101110;
20'b00101111110011101110: color_data = 12'b111011101110;
20'b00101111110011101111: color_data = 12'b111011101110;
20'b00101111110011110000: color_data = 12'b111011101110;
20'b00101111110011110001: color_data = 12'b111011101110;
20'b00101111110011110010: color_data = 12'b111011101110;
20'b00101111110011110011: color_data = 12'b111011101110;
20'b00101111110011110100: color_data = 12'b111011101110;
20'b00101111110011110101: color_data = 12'b111011101110;
20'b00101111110011110110: color_data = 12'b111011101110;
20'b00101111110011110111: color_data = 12'b111011101110;
20'b00101111110011111001: color_data = 12'b111011101110;
20'b00101111110011111010: color_data = 12'b111011101110;
20'b00101111110011111011: color_data = 12'b111011101110;
20'b00101111110011111100: color_data = 12'b111011101110;
20'b00101111110011111101: color_data = 12'b111011101110;
20'b00101111110011111110: color_data = 12'b111011101110;
20'b00101111110011111111: color_data = 12'b111011101110;
20'b00101111110100000000: color_data = 12'b111011101110;
20'b00101111110100000001: color_data = 12'b111011101110;
20'b00101111110100000010: color_data = 12'b111011101110;
20'b00101111110100100101: color_data = 12'b111011101110;
20'b00101111110100100110: color_data = 12'b111011101110;
20'b00101111110100100111: color_data = 12'b111011101110;
20'b00101111110100101000: color_data = 12'b111011101110;
20'b00101111110100101001: color_data = 12'b111011101110;
20'b00101111110100101010: color_data = 12'b111011101110;
20'b00101111110100101011: color_data = 12'b111011101110;
20'b00101111110100101100: color_data = 12'b111011101110;
20'b00101111110100101101: color_data = 12'b111011101110;
20'b00101111110100101110: color_data = 12'b111011101110;
20'b00101111110100110000: color_data = 12'b111011101110;
20'b00101111110100110001: color_data = 12'b111011101110;
20'b00101111110100110010: color_data = 12'b111011101110;
20'b00101111110100110011: color_data = 12'b111011101110;
20'b00101111110100110100: color_data = 12'b111011101110;
20'b00101111110100110101: color_data = 12'b111011101110;
20'b00101111110100110110: color_data = 12'b111011101110;
20'b00101111110100110111: color_data = 12'b111011101110;
20'b00101111110100111000: color_data = 12'b111011101110;
20'b00101111110100111001: color_data = 12'b111011101110;
20'b00101111110101000110: color_data = 12'b111011101110;
20'b00101111110101000111: color_data = 12'b111011101110;
20'b00101111110101001000: color_data = 12'b111011101110;
20'b00101111110101001001: color_data = 12'b111011101110;
20'b00101111110101001010: color_data = 12'b111011101110;
20'b00101111110101001011: color_data = 12'b111011101110;
20'b00101111110101001100: color_data = 12'b111011101110;
20'b00101111110101001101: color_data = 12'b111011101110;
20'b00101111110101001110: color_data = 12'b111011101110;
20'b00101111110101001111: color_data = 12'b111011101110;
20'b00101111110101010001: color_data = 12'b111011101110;
20'b00101111110101010010: color_data = 12'b111011101110;
20'b00101111110101010011: color_data = 12'b111011101110;
20'b00101111110101010100: color_data = 12'b111011101110;
20'b00101111110101010101: color_data = 12'b111011101110;
20'b00101111110101010110: color_data = 12'b111011101110;
20'b00101111110101010111: color_data = 12'b111011101110;
20'b00101111110101011000: color_data = 12'b111011101110;
20'b00101111110101011001: color_data = 12'b111011101110;
20'b00101111110101011010: color_data = 12'b111011101110;
20'b00101111110101111101: color_data = 12'b111011101110;
20'b00101111110101111110: color_data = 12'b111011101110;
20'b00101111110101111111: color_data = 12'b111011101110;
20'b00101111110110000000: color_data = 12'b111011101110;
20'b00101111110110000001: color_data = 12'b111011101110;
20'b00101111110110000010: color_data = 12'b111011101110;
20'b00101111110110000011: color_data = 12'b111011101110;
20'b00101111110110000100: color_data = 12'b111011101110;
20'b00101111110110000101: color_data = 12'b111011101110;
20'b00101111110110000110: color_data = 12'b111011101110;
20'b00101111110110001000: color_data = 12'b111011101110;
20'b00101111110110001001: color_data = 12'b111011101110;
20'b00101111110110001010: color_data = 12'b111011101110;
20'b00101111110110001011: color_data = 12'b111011101110;
20'b00101111110110001100: color_data = 12'b111011101110;
20'b00101111110110001101: color_data = 12'b111011101110;
20'b00101111110110001110: color_data = 12'b111011101110;
20'b00101111110110001111: color_data = 12'b111011101110;
20'b00101111110110010000: color_data = 12'b111011101110;
20'b00101111110110010001: color_data = 12'b111011101110;
20'b00101111110110011110: color_data = 12'b111011101110;
20'b00101111110110011111: color_data = 12'b111011101110;
20'b00101111110110100000: color_data = 12'b111011101110;
20'b00101111110110100001: color_data = 12'b111011101110;
20'b00101111110110100010: color_data = 12'b111011101110;
20'b00101111110110100011: color_data = 12'b111011101110;
20'b00101111110110100100: color_data = 12'b111011101110;
20'b00101111110110100101: color_data = 12'b111011101110;
20'b00101111110110100110: color_data = 12'b111011101110;
20'b00101111110110100111: color_data = 12'b111011101110;
20'b00101111110110101001: color_data = 12'b111011101110;
20'b00101111110110101010: color_data = 12'b111011101110;
20'b00101111110110101011: color_data = 12'b111011101110;
20'b00101111110110101100: color_data = 12'b111011101110;
20'b00101111110110101101: color_data = 12'b111011101110;
20'b00101111110110101110: color_data = 12'b111011101110;
20'b00101111110110101111: color_data = 12'b111011101110;
20'b00101111110110110000: color_data = 12'b111011101110;
20'b00101111110110110001: color_data = 12'b111011101110;
20'b00101111110110110010: color_data = 12'b111011101110;
20'b00101111110110110100: color_data = 12'b111011101110;
20'b00101111110110110101: color_data = 12'b111011101110;
20'b00101111110110110110: color_data = 12'b111011101110;
20'b00101111110110110111: color_data = 12'b111011101110;
20'b00101111110110111000: color_data = 12'b111011101110;
20'b00101111110110111001: color_data = 12'b111011101110;
20'b00101111110110111010: color_data = 12'b111011101110;
20'b00101111110110111011: color_data = 12'b111011101110;
20'b00101111110110111100: color_data = 12'b111011101110;
20'b00101111110110111101: color_data = 12'b111011101110;
20'b00101111110110111111: color_data = 12'b111011101110;
20'b00101111110111000000: color_data = 12'b111011101110;
20'b00101111110111000001: color_data = 12'b111011101110;
20'b00101111110111000010: color_data = 12'b111011101110;
20'b00101111110111000011: color_data = 12'b111011101110;
20'b00101111110111000100: color_data = 12'b111011101110;
20'b00101111110111000101: color_data = 12'b111011101110;
20'b00101111110111000110: color_data = 12'b111011101110;
20'b00101111110111000111: color_data = 12'b111011101110;
20'b00101111110111001000: color_data = 12'b111011101110;
20'b00101111110111001010: color_data = 12'b111011101110;
20'b00101111110111001011: color_data = 12'b111011101110;
20'b00101111110111001100: color_data = 12'b111011101110;
20'b00101111110111001101: color_data = 12'b111011101110;
20'b00101111110111001110: color_data = 12'b111011101110;
20'b00101111110111001111: color_data = 12'b111011101110;
20'b00101111110111010000: color_data = 12'b111011101110;
20'b00101111110111010001: color_data = 12'b111011101110;
20'b00101111110111010010: color_data = 12'b111011101110;
20'b00101111110111010011: color_data = 12'b111011101110;
20'b00101111110111010101: color_data = 12'b111011101110;
20'b00101111110111010110: color_data = 12'b111011101110;
20'b00101111110111010111: color_data = 12'b111011101110;
20'b00101111110111011000: color_data = 12'b111011101110;
20'b00101111110111011001: color_data = 12'b111011101110;
20'b00101111110111011010: color_data = 12'b111011101110;
20'b00101111110111011011: color_data = 12'b111011101110;
20'b00101111110111011100: color_data = 12'b111011101110;
20'b00101111110111011101: color_data = 12'b111011101110;
20'b00101111110111011110: color_data = 12'b111011101110;
20'b00101111110111100000: color_data = 12'b111011101110;
20'b00101111110111100001: color_data = 12'b111011101110;
20'b00101111110111100010: color_data = 12'b111011101110;
20'b00101111110111100011: color_data = 12'b111011101110;
20'b00101111110111100100: color_data = 12'b111011101110;
20'b00101111110111100101: color_data = 12'b111011101110;
20'b00101111110111100110: color_data = 12'b111011101110;
20'b00101111110111100111: color_data = 12'b111011101110;
20'b00101111110111101000: color_data = 12'b111011101110;
20'b00101111110111101001: color_data = 12'b111011101110;
20'b00110000000010100001: color_data = 12'b111011101110;
20'b00110000000010100010: color_data = 12'b111011101110;
20'b00110000000010100011: color_data = 12'b111011101110;
20'b00110000000010100100: color_data = 12'b111011101110;
20'b00110000000010100101: color_data = 12'b111011101110;
20'b00110000000010100110: color_data = 12'b111011101110;
20'b00110000000010100111: color_data = 12'b111011101110;
20'b00110000000010101000: color_data = 12'b111011101110;
20'b00110000000010101001: color_data = 12'b111011101110;
20'b00110000000010101010: color_data = 12'b111011101110;
20'b00110000000010101100: color_data = 12'b111011101110;
20'b00110000000010101101: color_data = 12'b111011101110;
20'b00110000000010101110: color_data = 12'b111011101110;
20'b00110000000010101111: color_data = 12'b111011101110;
20'b00110000000010110000: color_data = 12'b111011101110;
20'b00110000000010110001: color_data = 12'b111011101110;
20'b00110000000010110010: color_data = 12'b111011101110;
20'b00110000000010110011: color_data = 12'b111011101110;
20'b00110000000010110100: color_data = 12'b111011101110;
20'b00110000000010110101: color_data = 12'b111011101110;
20'b00110000000010110111: color_data = 12'b111011101110;
20'b00110000000010111000: color_data = 12'b111011101110;
20'b00110000000010111001: color_data = 12'b111011101110;
20'b00110000000010111010: color_data = 12'b111011101110;
20'b00110000000010111011: color_data = 12'b111011101110;
20'b00110000000010111100: color_data = 12'b111011101110;
20'b00110000000010111101: color_data = 12'b111011101110;
20'b00110000000010111110: color_data = 12'b111011101110;
20'b00110000000010111111: color_data = 12'b111011101110;
20'b00110000000011000000: color_data = 12'b111011101110;
20'b00110000000011000010: color_data = 12'b111011101110;
20'b00110000000011000011: color_data = 12'b111011101110;
20'b00110000000011000100: color_data = 12'b111011101110;
20'b00110000000011000101: color_data = 12'b111011101110;
20'b00110000000011000110: color_data = 12'b111011101110;
20'b00110000000011000111: color_data = 12'b111011101110;
20'b00110000000011001000: color_data = 12'b111011101110;
20'b00110000000011001001: color_data = 12'b111011101110;
20'b00110000000011001010: color_data = 12'b111011101110;
20'b00110000000011001011: color_data = 12'b111011101110;
20'b00110000000011001101: color_data = 12'b111011101110;
20'b00110000000011001110: color_data = 12'b111011101110;
20'b00110000000011001111: color_data = 12'b111011101110;
20'b00110000000011010000: color_data = 12'b111011101110;
20'b00110000000011010001: color_data = 12'b111011101110;
20'b00110000000011010010: color_data = 12'b111011101110;
20'b00110000000011010011: color_data = 12'b111011101110;
20'b00110000000011010100: color_data = 12'b111011101110;
20'b00110000000011010101: color_data = 12'b111011101110;
20'b00110000000011010110: color_data = 12'b111011101110;
20'b00110000000011101110: color_data = 12'b111011101110;
20'b00110000000011101111: color_data = 12'b111011101110;
20'b00110000000011110000: color_data = 12'b111011101110;
20'b00110000000011110001: color_data = 12'b111011101110;
20'b00110000000011110010: color_data = 12'b111011101110;
20'b00110000000011110011: color_data = 12'b111011101110;
20'b00110000000011110100: color_data = 12'b111011101110;
20'b00110000000011110101: color_data = 12'b111011101110;
20'b00110000000011110110: color_data = 12'b111011101110;
20'b00110000000011110111: color_data = 12'b111011101110;
20'b00110000000011111001: color_data = 12'b111011101110;
20'b00110000000011111010: color_data = 12'b111011101110;
20'b00110000000011111011: color_data = 12'b111011101110;
20'b00110000000011111100: color_data = 12'b111011101110;
20'b00110000000011111101: color_data = 12'b111011101110;
20'b00110000000011111110: color_data = 12'b111011101110;
20'b00110000000011111111: color_data = 12'b111011101110;
20'b00110000000100000000: color_data = 12'b111011101110;
20'b00110000000100000001: color_data = 12'b111011101110;
20'b00110000000100000010: color_data = 12'b111011101110;
20'b00110000000100100101: color_data = 12'b111011101110;
20'b00110000000100100110: color_data = 12'b111011101110;
20'b00110000000100100111: color_data = 12'b111011101110;
20'b00110000000100101000: color_data = 12'b111011101110;
20'b00110000000100101001: color_data = 12'b111011101110;
20'b00110000000100101010: color_data = 12'b111011101110;
20'b00110000000100101011: color_data = 12'b111011101110;
20'b00110000000100101100: color_data = 12'b111011101110;
20'b00110000000100101101: color_data = 12'b111011101110;
20'b00110000000100101110: color_data = 12'b111011101110;
20'b00110000000100110000: color_data = 12'b111011101110;
20'b00110000000100110001: color_data = 12'b111011101110;
20'b00110000000100110010: color_data = 12'b111011101110;
20'b00110000000100110011: color_data = 12'b111011101110;
20'b00110000000100110100: color_data = 12'b111011101110;
20'b00110000000100110101: color_data = 12'b111011101110;
20'b00110000000100110110: color_data = 12'b111011101110;
20'b00110000000100110111: color_data = 12'b111011101110;
20'b00110000000100111000: color_data = 12'b111011101110;
20'b00110000000100111001: color_data = 12'b111011101110;
20'b00110000000101000110: color_data = 12'b111011101110;
20'b00110000000101000111: color_data = 12'b111011101110;
20'b00110000000101001000: color_data = 12'b111011101110;
20'b00110000000101001001: color_data = 12'b111011101110;
20'b00110000000101001010: color_data = 12'b111011101110;
20'b00110000000101001011: color_data = 12'b111011101110;
20'b00110000000101001100: color_data = 12'b111011101110;
20'b00110000000101001101: color_data = 12'b111011101110;
20'b00110000000101001110: color_data = 12'b111011101110;
20'b00110000000101001111: color_data = 12'b111011101110;
20'b00110000000101010001: color_data = 12'b111011101110;
20'b00110000000101010010: color_data = 12'b111011101110;
20'b00110000000101010011: color_data = 12'b111011101110;
20'b00110000000101010100: color_data = 12'b111011101110;
20'b00110000000101010101: color_data = 12'b111011101110;
20'b00110000000101010110: color_data = 12'b111011101110;
20'b00110000000101010111: color_data = 12'b111011101110;
20'b00110000000101011000: color_data = 12'b111011101110;
20'b00110000000101011001: color_data = 12'b111011101110;
20'b00110000000101011010: color_data = 12'b111011101110;
20'b00110000000101111101: color_data = 12'b111011101110;
20'b00110000000101111110: color_data = 12'b111011101110;
20'b00110000000101111111: color_data = 12'b111011101110;
20'b00110000000110000000: color_data = 12'b111011101110;
20'b00110000000110000001: color_data = 12'b111011101110;
20'b00110000000110000010: color_data = 12'b111011101110;
20'b00110000000110000011: color_data = 12'b111011101110;
20'b00110000000110000100: color_data = 12'b111011101110;
20'b00110000000110000101: color_data = 12'b111011101110;
20'b00110000000110000110: color_data = 12'b111011101110;
20'b00110000000110001000: color_data = 12'b111011101110;
20'b00110000000110001001: color_data = 12'b111011101110;
20'b00110000000110001010: color_data = 12'b111011101110;
20'b00110000000110001011: color_data = 12'b111011101110;
20'b00110000000110001100: color_data = 12'b111011101110;
20'b00110000000110001101: color_data = 12'b111011101110;
20'b00110000000110001110: color_data = 12'b111011101110;
20'b00110000000110001111: color_data = 12'b111011101110;
20'b00110000000110010000: color_data = 12'b111011101110;
20'b00110000000110010001: color_data = 12'b111011101110;
20'b00110000000110011110: color_data = 12'b111011101110;
20'b00110000000110011111: color_data = 12'b111011101110;
20'b00110000000110100000: color_data = 12'b111011101110;
20'b00110000000110100001: color_data = 12'b111011101110;
20'b00110000000110100010: color_data = 12'b111011101110;
20'b00110000000110100011: color_data = 12'b111011101110;
20'b00110000000110100100: color_data = 12'b111011101110;
20'b00110000000110100101: color_data = 12'b111011101110;
20'b00110000000110100110: color_data = 12'b111011101110;
20'b00110000000110100111: color_data = 12'b111011101110;
20'b00110000000110101001: color_data = 12'b111011101110;
20'b00110000000110101010: color_data = 12'b111011101110;
20'b00110000000110101011: color_data = 12'b111011101110;
20'b00110000000110101100: color_data = 12'b111011101110;
20'b00110000000110101101: color_data = 12'b111011101110;
20'b00110000000110101110: color_data = 12'b111011101110;
20'b00110000000110101111: color_data = 12'b111011101110;
20'b00110000000110110000: color_data = 12'b111011101110;
20'b00110000000110110001: color_data = 12'b111011101110;
20'b00110000000110110010: color_data = 12'b111011101110;
20'b00110000000110110100: color_data = 12'b111011101110;
20'b00110000000110110101: color_data = 12'b111011101110;
20'b00110000000110110110: color_data = 12'b111011101110;
20'b00110000000110110111: color_data = 12'b111011101110;
20'b00110000000110111000: color_data = 12'b111011101110;
20'b00110000000110111001: color_data = 12'b111011101110;
20'b00110000000110111010: color_data = 12'b111011101110;
20'b00110000000110111011: color_data = 12'b111011101110;
20'b00110000000110111100: color_data = 12'b111011101110;
20'b00110000000110111101: color_data = 12'b111011101110;
20'b00110000000110111111: color_data = 12'b111011101110;
20'b00110000000111000000: color_data = 12'b111011101110;
20'b00110000000111000001: color_data = 12'b111011101110;
20'b00110000000111000010: color_data = 12'b111011101110;
20'b00110000000111000011: color_data = 12'b111011101110;
20'b00110000000111000100: color_data = 12'b111011101110;
20'b00110000000111000101: color_data = 12'b111011101110;
20'b00110000000111000110: color_data = 12'b111011101110;
20'b00110000000111000111: color_data = 12'b111011101110;
20'b00110000000111001000: color_data = 12'b111011101110;
20'b00110000000111001010: color_data = 12'b111011101110;
20'b00110000000111001011: color_data = 12'b111011101110;
20'b00110000000111001100: color_data = 12'b111011101110;
20'b00110000000111001101: color_data = 12'b111011101110;
20'b00110000000111001110: color_data = 12'b111011101110;
20'b00110000000111001111: color_data = 12'b111011101110;
20'b00110000000111010000: color_data = 12'b111011101110;
20'b00110000000111010001: color_data = 12'b111011101110;
20'b00110000000111010010: color_data = 12'b111011101110;
20'b00110000000111010011: color_data = 12'b111011101110;
20'b00110000000111010101: color_data = 12'b111011101110;
20'b00110000000111010110: color_data = 12'b111011101110;
20'b00110000000111010111: color_data = 12'b111011101110;
20'b00110000000111011000: color_data = 12'b111011101110;
20'b00110000000111011001: color_data = 12'b111011101110;
20'b00110000000111011010: color_data = 12'b111011101110;
20'b00110000000111011011: color_data = 12'b111011101110;
20'b00110000000111011100: color_data = 12'b111011101110;
20'b00110000000111011101: color_data = 12'b111011101110;
20'b00110000000111011110: color_data = 12'b111011101110;
20'b00110000000111100000: color_data = 12'b111011101110;
20'b00110000000111100001: color_data = 12'b111011101110;
20'b00110000000111100010: color_data = 12'b111011101110;
20'b00110000000111100011: color_data = 12'b111011101110;
20'b00110000000111100100: color_data = 12'b111011101110;
20'b00110000000111100101: color_data = 12'b111011101110;
20'b00110000000111100110: color_data = 12'b111011101110;
20'b00110000000111100111: color_data = 12'b111011101110;
20'b00110000000111101000: color_data = 12'b111011101110;
20'b00110000000111101001: color_data = 12'b111011101110;
20'b00110000010010100001: color_data = 12'b111011101110;
20'b00110000010010100010: color_data = 12'b111011101110;
20'b00110000010010100011: color_data = 12'b111011101110;
20'b00110000010010100100: color_data = 12'b111011101110;
20'b00110000010010100101: color_data = 12'b111011101110;
20'b00110000010010100110: color_data = 12'b111011101110;
20'b00110000010010100111: color_data = 12'b111011101110;
20'b00110000010010101000: color_data = 12'b111011101110;
20'b00110000010010101001: color_data = 12'b111011101110;
20'b00110000010010101010: color_data = 12'b111011101110;
20'b00110000010010101100: color_data = 12'b111011101110;
20'b00110000010010101101: color_data = 12'b111011101110;
20'b00110000010010101110: color_data = 12'b111011101110;
20'b00110000010010101111: color_data = 12'b111011101110;
20'b00110000010010110000: color_data = 12'b111011101110;
20'b00110000010010110001: color_data = 12'b111011101110;
20'b00110000010010110010: color_data = 12'b111011101110;
20'b00110000010010110011: color_data = 12'b111011101110;
20'b00110000010010110100: color_data = 12'b111011101110;
20'b00110000010010110101: color_data = 12'b111011101110;
20'b00110000010010110111: color_data = 12'b111011101110;
20'b00110000010010111000: color_data = 12'b111011101110;
20'b00110000010010111001: color_data = 12'b111011101110;
20'b00110000010010111010: color_data = 12'b111011101110;
20'b00110000010010111011: color_data = 12'b111011101110;
20'b00110000010010111100: color_data = 12'b111011101110;
20'b00110000010010111101: color_data = 12'b111011101110;
20'b00110000010010111110: color_data = 12'b111011101110;
20'b00110000010010111111: color_data = 12'b111011101110;
20'b00110000010011000000: color_data = 12'b111011101110;
20'b00110000010011000010: color_data = 12'b111011101110;
20'b00110000010011000011: color_data = 12'b111011101110;
20'b00110000010011000100: color_data = 12'b111011101110;
20'b00110000010011000101: color_data = 12'b111011101110;
20'b00110000010011000110: color_data = 12'b111011101110;
20'b00110000010011000111: color_data = 12'b111011101110;
20'b00110000010011001000: color_data = 12'b111011101110;
20'b00110000010011001001: color_data = 12'b111011101110;
20'b00110000010011001010: color_data = 12'b111011101110;
20'b00110000010011001011: color_data = 12'b111011101110;
20'b00110000010011001101: color_data = 12'b111011101110;
20'b00110000010011001110: color_data = 12'b111011101110;
20'b00110000010011001111: color_data = 12'b111011101110;
20'b00110000010011010000: color_data = 12'b111011101110;
20'b00110000010011010001: color_data = 12'b111011101110;
20'b00110000010011010010: color_data = 12'b111011101110;
20'b00110000010011010011: color_data = 12'b111011101110;
20'b00110000010011010100: color_data = 12'b111011101110;
20'b00110000010011010101: color_data = 12'b111011101110;
20'b00110000010011010110: color_data = 12'b111011101110;
20'b00110000010011101110: color_data = 12'b111011101110;
20'b00110000010011101111: color_data = 12'b111011101110;
20'b00110000010011110000: color_data = 12'b111011101110;
20'b00110000010011110001: color_data = 12'b111011101110;
20'b00110000010011110010: color_data = 12'b111011101110;
20'b00110000010011110011: color_data = 12'b111011101110;
20'b00110000010011110100: color_data = 12'b111011101110;
20'b00110000010011110101: color_data = 12'b111011101110;
20'b00110000010011110110: color_data = 12'b111011101110;
20'b00110000010011110111: color_data = 12'b111011101110;
20'b00110000010011111001: color_data = 12'b111011101110;
20'b00110000010011111010: color_data = 12'b111011101110;
20'b00110000010011111011: color_data = 12'b111011101110;
20'b00110000010011111100: color_data = 12'b111011101110;
20'b00110000010011111101: color_data = 12'b111011101110;
20'b00110000010011111110: color_data = 12'b111011101110;
20'b00110000010011111111: color_data = 12'b111011101110;
20'b00110000010100000000: color_data = 12'b111011101110;
20'b00110000010100000001: color_data = 12'b111011101110;
20'b00110000010100000010: color_data = 12'b111011101110;
20'b00110000010100100101: color_data = 12'b111011101110;
20'b00110000010100100110: color_data = 12'b111011101110;
20'b00110000010100100111: color_data = 12'b111011101110;
20'b00110000010100101000: color_data = 12'b111011101110;
20'b00110000010100101001: color_data = 12'b111011101110;
20'b00110000010100101010: color_data = 12'b111011101110;
20'b00110000010100101011: color_data = 12'b111011101110;
20'b00110000010100101100: color_data = 12'b111011101110;
20'b00110000010100101101: color_data = 12'b111011101110;
20'b00110000010100101110: color_data = 12'b111011101110;
20'b00110000010100110000: color_data = 12'b111011101110;
20'b00110000010100110001: color_data = 12'b111011101110;
20'b00110000010100110010: color_data = 12'b111011101110;
20'b00110000010100110011: color_data = 12'b111011101110;
20'b00110000010100110100: color_data = 12'b111011101110;
20'b00110000010100110101: color_data = 12'b111011101110;
20'b00110000010100110110: color_data = 12'b111011101110;
20'b00110000010100110111: color_data = 12'b111011101110;
20'b00110000010100111000: color_data = 12'b111011101110;
20'b00110000010100111001: color_data = 12'b111011101110;
20'b00110000010101000110: color_data = 12'b111011101110;
20'b00110000010101000111: color_data = 12'b111011101110;
20'b00110000010101001000: color_data = 12'b111011101110;
20'b00110000010101001001: color_data = 12'b111011101110;
20'b00110000010101001010: color_data = 12'b111011101110;
20'b00110000010101001011: color_data = 12'b111011101110;
20'b00110000010101001100: color_data = 12'b111011101110;
20'b00110000010101001101: color_data = 12'b111011101110;
20'b00110000010101001110: color_data = 12'b111011101110;
20'b00110000010101001111: color_data = 12'b111011101110;
20'b00110000010101010001: color_data = 12'b111011101110;
20'b00110000010101010010: color_data = 12'b111011101110;
20'b00110000010101010011: color_data = 12'b111011101110;
20'b00110000010101010100: color_data = 12'b111011101110;
20'b00110000010101010101: color_data = 12'b111011101110;
20'b00110000010101010110: color_data = 12'b111011101110;
20'b00110000010101010111: color_data = 12'b111011101110;
20'b00110000010101011000: color_data = 12'b111011101110;
20'b00110000010101011001: color_data = 12'b111011101110;
20'b00110000010101011010: color_data = 12'b111011101110;
20'b00110000010101111101: color_data = 12'b111011101110;
20'b00110000010101111110: color_data = 12'b111011101110;
20'b00110000010101111111: color_data = 12'b111011101110;
20'b00110000010110000000: color_data = 12'b111011101110;
20'b00110000010110000001: color_data = 12'b111011101110;
20'b00110000010110000010: color_data = 12'b111011101110;
20'b00110000010110000011: color_data = 12'b111011101110;
20'b00110000010110000100: color_data = 12'b111011101110;
20'b00110000010110000101: color_data = 12'b111011101110;
20'b00110000010110000110: color_data = 12'b111011101110;
20'b00110000010110001000: color_data = 12'b111011101110;
20'b00110000010110001001: color_data = 12'b111011101110;
20'b00110000010110001010: color_data = 12'b111011101110;
20'b00110000010110001011: color_data = 12'b111011101110;
20'b00110000010110001100: color_data = 12'b111011101110;
20'b00110000010110001101: color_data = 12'b111011101110;
20'b00110000010110001110: color_data = 12'b111011101110;
20'b00110000010110001111: color_data = 12'b111011101110;
20'b00110000010110010000: color_data = 12'b111011101110;
20'b00110000010110010001: color_data = 12'b111011101110;
20'b00110000010110011110: color_data = 12'b111011101110;
20'b00110000010110011111: color_data = 12'b111011101110;
20'b00110000010110100000: color_data = 12'b111011101110;
20'b00110000010110100001: color_data = 12'b111011101110;
20'b00110000010110100010: color_data = 12'b111011101110;
20'b00110000010110100011: color_data = 12'b111011101110;
20'b00110000010110100100: color_data = 12'b111011101110;
20'b00110000010110100101: color_data = 12'b111011101110;
20'b00110000010110100110: color_data = 12'b111011101110;
20'b00110000010110100111: color_data = 12'b111011101110;
20'b00110000010110101001: color_data = 12'b111011101110;
20'b00110000010110101010: color_data = 12'b111011101110;
20'b00110000010110101011: color_data = 12'b111011101110;
20'b00110000010110101100: color_data = 12'b111011101110;
20'b00110000010110101101: color_data = 12'b111011101110;
20'b00110000010110101110: color_data = 12'b111011101110;
20'b00110000010110101111: color_data = 12'b111011101110;
20'b00110000010110110000: color_data = 12'b111011101110;
20'b00110000010110110001: color_data = 12'b111011101110;
20'b00110000010110110010: color_data = 12'b111011101110;
20'b00110000010110110100: color_data = 12'b111011101110;
20'b00110000010110110101: color_data = 12'b111011101110;
20'b00110000010110110110: color_data = 12'b111011101110;
20'b00110000010110110111: color_data = 12'b111011101110;
20'b00110000010110111000: color_data = 12'b111011101110;
20'b00110000010110111001: color_data = 12'b111011101110;
20'b00110000010110111010: color_data = 12'b111011101110;
20'b00110000010110111011: color_data = 12'b111011101110;
20'b00110000010110111100: color_data = 12'b111011101110;
20'b00110000010110111101: color_data = 12'b111011101110;
20'b00110000010110111111: color_data = 12'b111011101110;
20'b00110000010111000000: color_data = 12'b111011101110;
20'b00110000010111000001: color_data = 12'b111011101110;
20'b00110000010111000010: color_data = 12'b111011101110;
20'b00110000010111000011: color_data = 12'b111011101110;
20'b00110000010111000100: color_data = 12'b111011101110;
20'b00110000010111000101: color_data = 12'b111011101110;
20'b00110000010111000110: color_data = 12'b111011101110;
20'b00110000010111000111: color_data = 12'b111011101110;
20'b00110000010111001000: color_data = 12'b111011101110;
20'b00110000010111001010: color_data = 12'b111011101110;
20'b00110000010111001011: color_data = 12'b111011101110;
20'b00110000010111001100: color_data = 12'b111011101110;
20'b00110000010111001101: color_data = 12'b111011101110;
20'b00110000010111001110: color_data = 12'b111011101110;
20'b00110000010111001111: color_data = 12'b111011101110;
20'b00110000010111010000: color_data = 12'b111011101110;
20'b00110000010111010001: color_data = 12'b111011101110;
20'b00110000010111010010: color_data = 12'b111011101110;
20'b00110000010111010011: color_data = 12'b111011101110;
20'b00110000010111010101: color_data = 12'b111011101110;
20'b00110000010111010110: color_data = 12'b111011101110;
20'b00110000010111010111: color_data = 12'b111011101110;
20'b00110000010111011000: color_data = 12'b111011101110;
20'b00110000010111011001: color_data = 12'b111011101110;
20'b00110000010111011010: color_data = 12'b111011101110;
20'b00110000010111011011: color_data = 12'b111011101110;
20'b00110000010111011100: color_data = 12'b111011101110;
20'b00110000010111011101: color_data = 12'b111011101110;
20'b00110000010111011110: color_data = 12'b111011101110;
20'b00110000010111100000: color_data = 12'b111011101110;
20'b00110000010111100001: color_data = 12'b111011101110;
20'b00110000010111100010: color_data = 12'b111011101110;
20'b00110000010111100011: color_data = 12'b111011101110;
20'b00110000010111100100: color_data = 12'b111011101110;
20'b00110000010111100101: color_data = 12'b111011101110;
20'b00110000010111100110: color_data = 12'b111011101110;
20'b00110000010111100111: color_data = 12'b111011101110;
20'b00110000010111101000: color_data = 12'b111011101110;
20'b00110000010111101001: color_data = 12'b111011101110;
20'b00110000100010100001: color_data = 12'b111011101110;
20'b00110000100010100010: color_data = 12'b111011101110;
20'b00110000100010100011: color_data = 12'b111011101110;
20'b00110000100010100100: color_data = 12'b111011101110;
20'b00110000100010100101: color_data = 12'b111011101110;
20'b00110000100010100110: color_data = 12'b111011101110;
20'b00110000100010100111: color_data = 12'b111011101110;
20'b00110000100010101000: color_data = 12'b111011101110;
20'b00110000100010101001: color_data = 12'b111011101110;
20'b00110000100010101010: color_data = 12'b111011101110;
20'b00110000100010101100: color_data = 12'b111011101110;
20'b00110000100010101101: color_data = 12'b111011101110;
20'b00110000100010101110: color_data = 12'b111011101110;
20'b00110000100010101111: color_data = 12'b111011101110;
20'b00110000100010110000: color_data = 12'b111011101110;
20'b00110000100010110001: color_data = 12'b111011101110;
20'b00110000100010110010: color_data = 12'b111011101110;
20'b00110000100010110011: color_data = 12'b111011101110;
20'b00110000100010110100: color_data = 12'b111011101110;
20'b00110000100010110101: color_data = 12'b111011101110;
20'b00110000100010110111: color_data = 12'b111011101110;
20'b00110000100010111000: color_data = 12'b111011101110;
20'b00110000100010111001: color_data = 12'b111011101110;
20'b00110000100010111010: color_data = 12'b111011101110;
20'b00110000100010111011: color_data = 12'b111011101110;
20'b00110000100010111100: color_data = 12'b111011101110;
20'b00110000100010111101: color_data = 12'b111011101110;
20'b00110000100010111110: color_data = 12'b111011101110;
20'b00110000100010111111: color_data = 12'b111011101110;
20'b00110000100011000000: color_data = 12'b111011101110;
20'b00110000100011000010: color_data = 12'b111011101110;
20'b00110000100011000011: color_data = 12'b111011101110;
20'b00110000100011000100: color_data = 12'b111011101110;
20'b00110000100011000101: color_data = 12'b111011101110;
20'b00110000100011000110: color_data = 12'b111011101110;
20'b00110000100011000111: color_data = 12'b111011101110;
20'b00110000100011001000: color_data = 12'b111011101110;
20'b00110000100011001001: color_data = 12'b111011101110;
20'b00110000100011001010: color_data = 12'b111011101110;
20'b00110000100011001011: color_data = 12'b111011101110;
20'b00110000100011001101: color_data = 12'b111011101110;
20'b00110000100011001110: color_data = 12'b111011101110;
20'b00110000100011001111: color_data = 12'b111011101110;
20'b00110000100011010000: color_data = 12'b111011101110;
20'b00110000100011010001: color_data = 12'b111011101110;
20'b00110000100011010010: color_data = 12'b111011101110;
20'b00110000100011010011: color_data = 12'b111011101110;
20'b00110000100011010100: color_data = 12'b111011101110;
20'b00110000100011010101: color_data = 12'b111011101110;
20'b00110000100011010110: color_data = 12'b111011101110;
20'b00110000100011101110: color_data = 12'b111011101110;
20'b00110000100011101111: color_data = 12'b111011101110;
20'b00110000100011110000: color_data = 12'b111011101110;
20'b00110000100011110001: color_data = 12'b111011101110;
20'b00110000100011110010: color_data = 12'b111011101110;
20'b00110000100011110011: color_data = 12'b111011101110;
20'b00110000100011110100: color_data = 12'b111011101110;
20'b00110000100011110101: color_data = 12'b111011101110;
20'b00110000100011110110: color_data = 12'b111011101110;
20'b00110000100011110111: color_data = 12'b111011101110;
20'b00110000100011111001: color_data = 12'b111011101110;
20'b00110000100011111010: color_data = 12'b111011101110;
20'b00110000100011111011: color_data = 12'b111011101110;
20'b00110000100011111100: color_data = 12'b111011101110;
20'b00110000100011111101: color_data = 12'b111011101110;
20'b00110000100011111110: color_data = 12'b111011101110;
20'b00110000100011111111: color_data = 12'b111011101110;
20'b00110000100100000000: color_data = 12'b111011101110;
20'b00110000100100000001: color_data = 12'b111011101110;
20'b00110000100100000010: color_data = 12'b111011101110;
20'b00110000100100100101: color_data = 12'b111011101110;
20'b00110000100100100110: color_data = 12'b111011101110;
20'b00110000100100100111: color_data = 12'b111011101110;
20'b00110000100100101000: color_data = 12'b111011101110;
20'b00110000100100101001: color_data = 12'b111011101110;
20'b00110000100100101010: color_data = 12'b111011101110;
20'b00110000100100101011: color_data = 12'b111011101110;
20'b00110000100100101100: color_data = 12'b111011101110;
20'b00110000100100101101: color_data = 12'b111011101110;
20'b00110000100100101110: color_data = 12'b111011101110;
20'b00110000100100110000: color_data = 12'b111011101110;
20'b00110000100100110001: color_data = 12'b111011101110;
20'b00110000100100110010: color_data = 12'b111011101110;
20'b00110000100100110011: color_data = 12'b111011101110;
20'b00110000100100110100: color_data = 12'b111011101110;
20'b00110000100100110101: color_data = 12'b111011101110;
20'b00110000100100110110: color_data = 12'b111011101110;
20'b00110000100100110111: color_data = 12'b111011101110;
20'b00110000100100111000: color_data = 12'b111011101110;
20'b00110000100100111001: color_data = 12'b111011101110;
20'b00110000100101000110: color_data = 12'b111011101110;
20'b00110000100101000111: color_data = 12'b111011101110;
20'b00110000100101001000: color_data = 12'b111011101110;
20'b00110000100101001001: color_data = 12'b111011101110;
20'b00110000100101001010: color_data = 12'b111011101110;
20'b00110000100101001011: color_data = 12'b111011101110;
20'b00110000100101001100: color_data = 12'b111011101110;
20'b00110000100101001101: color_data = 12'b111011101110;
20'b00110000100101001110: color_data = 12'b111011101110;
20'b00110000100101001111: color_data = 12'b111011101110;
20'b00110000100101010001: color_data = 12'b111011101110;
20'b00110000100101010010: color_data = 12'b111011101110;
20'b00110000100101010011: color_data = 12'b111011101110;
20'b00110000100101010100: color_data = 12'b111011101110;
20'b00110000100101010101: color_data = 12'b111011101110;
20'b00110000100101010110: color_data = 12'b111011101110;
20'b00110000100101010111: color_data = 12'b111011101110;
20'b00110000100101011000: color_data = 12'b111011101110;
20'b00110000100101011001: color_data = 12'b111011101110;
20'b00110000100101011010: color_data = 12'b111011101110;
20'b00110000100101111101: color_data = 12'b111011101110;
20'b00110000100101111110: color_data = 12'b111011101110;
20'b00110000100101111111: color_data = 12'b111011101110;
20'b00110000100110000000: color_data = 12'b111011101110;
20'b00110000100110000001: color_data = 12'b111011101110;
20'b00110000100110000010: color_data = 12'b111011101110;
20'b00110000100110000011: color_data = 12'b111011101110;
20'b00110000100110000100: color_data = 12'b111011101110;
20'b00110000100110000101: color_data = 12'b111011101110;
20'b00110000100110000110: color_data = 12'b111011101110;
20'b00110000100110001000: color_data = 12'b111011101110;
20'b00110000100110001001: color_data = 12'b111011101110;
20'b00110000100110001010: color_data = 12'b111011101110;
20'b00110000100110001011: color_data = 12'b111011101110;
20'b00110000100110001100: color_data = 12'b111011101110;
20'b00110000100110001101: color_data = 12'b111011101110;
20'b00110000100110001110: color_data = 12'b111011101110;
20'b00110000100110001111: color_data = 12'b111011101110;
20'b00110000100110010000: color_data = 12'b111011101110;
20'b00110000100110010001: color_data = 12'b111011101110;
20'b00110000100110011110: color_data = 12'b111011101110;
20'b00110000100110011111: color_data = 12'b111011101110;
20'b00110000100110100000: color_data = 12'b111011101110;
20'b00110000100110100001: color_data = 12'b111011101110;
20'b00110000100110100010: color_data = 12'b111011101110;
20'b00110000100110100011: color_data = 12'b111011101110;
20'b00110000100110100100: color_data = 12'b111011101110;
20'b00110000100110100101: color_data = 12'b111011101110;
20'b00110000100110100110: color_data = 12'b111011101110;
20'b00110000100110100111: color_data = 12'b111011101110;
20'b00110000100110101001: color_data = 12'b111011101110;
20'b00110000100110101010: color_data = 12'b111011101110;
20'b00110000100110101011: color_data = 12'b111011101110;
20'b00110000100110101100: color_data = 12'b111011101110;
20'b00110000100110101101: color_data = 12'b111011101110;
20'b00110000100110101110: color_data = 12'b111011101110;
20'b00110000100110101111: color_data = 12'b111011101110;
20'b00110000100110110000: color_data = 12'b111011101110;
20'b00110000100110110001: color_data = 12'b111011101110;
20'b00110000100110110010: color_data = 12'b111011101110;
20'b00110000100110110100: color_data = 12'b111011101110;
20'b00110000100110110101: color_data = 12'b111011101110;
20'b00110000100110110110: color_data = 12'b111011101110;
20'b00110000100110110111: color_data = 12'b111011101110;
20'b00110000100110111000: color_data = 12'b111011101110;
20'b00110000100110111001: color_data = 12'b111011101110;
20'b00110000100110111010: color_data = 12'b111011101110;
20'b00110000100110111011: color_data = 12'b111011101110;
20'b00110000100110111100: color_data = 12'b111011101110;
20'b00110000100110111101: color_data = 12'b111011101110;
20'b00110000100110111111: color_data = 12'b111011101110;
20'b00110000100111000000: color_data = 12'b111011101110;
20'b00110000100111000001: color_data = 12'b111011101110;
20'b00110000100111000010: color_data = 12'b111011101110;
20'b00110000100111000011: color_data = 12'b111011101110;
20'b00110000100111000100: color_data = 12'b111011101110;
20'b00110000100111000101: color_data = 12'b111011101110;
20'b00110000100111000110: color_data = 12'b111011101110;
20'b00110000100111000111: color_data = 12'b111011101110;
20'b00110000100111001000: color_data = 12'b111011101110;
20'b00110000100111001010: color_data = 12'b111011101110;
20'b00110000100111001011: color_data = 12'b111011101110;
20'b00110000100111001100: color_data = 12'b111011101110;
20'b00110000100111001101: color_data = 12'b111011101110;
20'b00110000100111001110: color_data = 12'b111011101110;
20'b00110000100111001111: color_data = 12'b111011101110;
20'b00110000100111010000: color_data = 12'b111011101110;
20'b00110000100111010001: color_data = 12'b111011101110;
20'b00110000100111010010: color_data = 12'b111011101110;
20'b00110000100111010011: color_data = 12'b111011101110;
20'b00110000100111010101: color_data = 12'b111011101110;
20'b00110000100111010110: color_data = 12'b111011101110;
20'b00110000100111010111: color_data = 12'b111011101110;
20'b00110000100111011000: color_data = 12'b111011101110;
20'b00110000100111011001: color_data = 12'b111011101110;
20'b00110000100111011010: color_data = 12'b111011101110;
20'b00110000100111011011: color_data = 12'b111011101110;
20'b00110000100111011100: color_data = 12'b111011101110;
20'b00110000100111011101: color_data = 12'b111011101110;
20'b00110000100111011110: color_data = 12'b111011101110;
20'b00110000100111100000: color_data = 12'b111011101110;
20'b00110000100111100001: color_data = 12'b111011101110;
20'b00110000100111100010: color_data = 12'b111011101110;
20'b00110000100111100011: color_data = 12'b111011101110;
20'b00110000100111100100: color_data = 12'b111011101110;
20'b00110000100111100101: color_data = 12'b111011101110;
20'b00110000100111100110: color_data = 12'b111011101110;
20'b00110000100111100111: color_data = 12'b111011101110;
20'b00110000100111101000: color_data = 12'b111011101110;
20'b00110000100111101001: color_data = 12'b111011101110;
20'b00110000110010100001: color_data = 12'b111011101110;
20'b00110000110010100010: color_data = 12'b111011101110;
20'b00110000110010100011: color_data = 12'b111011101110;
20'b00110000110010100100: color_data = 12'b111011101110;
20'b00110000110010100101: color_data = 12'b111011101110;
20'b00110000110010100110: color_data = 12'b111011101110;
20'b00110000110010100111: color_data = 12'b111011101110;
20'b00110000110010101000: color_data = 12'b111011101110;
20'b00110000110010101001: color_data = 12'b111011101110;
20'b00110000110010101010: color_data = 12'b111011101110;
20'b00110000110010101100: color_data = 12'b111011101110;
20'b00110000110010101101: color_data = 12'b111011101110;
20'b00110000110010101110: color_data = 12'b111011101110;
20'b00110000110010101111: color_data = 12'b111011101110;
20'b00110000110010110000: color_data = 12'b111011101110;
20'b00110000110010110001: color_data = 12'b111011101110;
20'b00110000110010110010: color_data = 12'b111011101110;
20'b00110000110010110011: color_data = 12'b111011101110;
20'b00110000110010110100: color_data = 12'b111011101110;
20'b00110000110010110101: color_data = 12'b111011101110;
20'b00110000110010110111: color_data = 12'b111011101110;
20'b00110000110010111000: color_data = 12'b111011101110;
20'b00110000110010111001: color_data = 12'b111011101110;
20'b00110000110010111010: color_data = 12'b111011101110;
20'b00110000110010111011: color_data = 12'b111011101110;
20'b00110000110010111100: color_data = 12'b111011101110;
20'b00110000110010111101: color_data = 12'b111011101110;
20'b00110000110010111110: color_data = 12'b111011101110;
20'b00110000110010111111: color_data = 12'b111011101110;
20'b00110000110011000000: color_data = 12'b111011101110;
20'b00110000110011000010: color_data = 12'b111011101110;
20'b00110000110011000011: color_data = 12'b111011101110;
20'b00110000110011000100: color_data = 12'b111011101110;
20'b00110000110011000101: color_data = 12'b111011101110;
20'b00110000110011000110: color_data = 12'b111011101110;
20'b00110000110011000111: color_data = 12'b111011101110;
20'b00110000110011001000: color_data = 12'b111011101110;
20'b00110000110011001001: color_data = 12'b111011101110;
20'b00110000110011001010: color_data = 12'b111011101110;
20'b00110000110011001011: color_data = 12'b111011101110;
20'b00110000110011001101: color_data = 12'b111011101110;
20'b00110000110011001110: color_data = 12'b111011101110;
20'b00110000110011001111: color_data = 12'b111011101110;
20'b00110000110011010000: color_data = 12'b111011101110;
20'b00110000110011010001: color_data = 12'b111011101110;
20'b00110000110011010010: color_data = 12'b111011101110;
20'b00110000110011010011: color_data = 12'b111011101110;
20'b00110000110011010100: color_data = 12'b111011101110;
20'b00110000110011010101: color_data = 12'b111011101110;
20'b00110000110011010110: color_data = 12'b111011101110;
20'b00110000110011101110: color_data = 12'b111011101110;
20'b00110000110011101111: color_data = 12'b111011101110;
20'b00110000110011110000: color_data = 12'b111011101110;
20'b00110000110011110001: color_data = 12'b111011101110;
20'b00110000110011110010: color_data = 12'b111011101110;
20'b00110000110011110011: color_data = 12'b111011101110;
20'b00110000110011110100: color_data = 12'b111011101110;
20'b00110000110011110101: color_data = 12'b111011101110;
20'b00110000110011110110: color_data = 12'b111011101110;
20'b00110000110011110111: color_data = 12'b111011101110;
20'b00110000110011111001: color_data = 12'b111011101110;
20'b00110000110011111010: color_data = 12'b111011101110;
20'b00110000110011111011: color_data = 12'b111011101110;
20'b00110000110011111100: color_data = 12'b111011101110;
20'b00110000110011111101: color_data = 12'b111011101110;
20'b00110000110011111110: color_data = 12'b111011101110;
20'b00110000110011111111: color_data = 12'b111011101110;
20'b00110000110100000000: color_data = 12'b111011101110;
20'b00110000110100000001: color_data = 12'b111011101110;
20'b00110000110100000010: color_data = 12'b111011101110;
20'b00110000110100100101: color_data = 12'b111011101110;
20'b00110000110100100110: color_data = 12'b111011101110;
20'b00110000110100100111: color_data = 12'b111011101110;
20'b00110000110100101000: color_data = 12'b111011101110;
20'b00110000110100101001: color_data = 12'b111011101110;
20'b00110000110100101010: color_data = 12'b111011101110;
20'b00110000110100101011: color_data = 12'b111011101110;
20'b00110000110100101100: color_data = 12'b111011101110;
20'b00110000110100101101: color_data = 12'b111011101110;
20'b00110000110100101110: color_data = 12'b111011101110;
20'b00110000110100110000: color_data = 12'b111011101110;
20'b00110000110100110001: color_data = 12'b111011101110;
20'b00110000110100110010: color_data = 12'b111011101110;
20'b00110000110100110011: color_data = 12'b111011101110;
20'b00110000110100110100: color_data = 12'b111011101110;
20'b00110000110100110101: color_data = 12'b111011101110;
20'b00110000110100110110: color_data = 12'b111011101110;
20'b00110000110100110111: color_data = 12'b111011101110;
20'b00110000110100111000: color_data = 12'b111011101110;
20'b00110000110100111001: color_data = 12'b111011101110;
20'b00110000110101000110: color_data = 12'b111011101110;
20'b00110000110101000111: color_data = 12'b111011101110;
20'b00110000110101001000: color_data = 12'b111011101110;
20'b00110000110101001001: color_data = 12'b111011101110;
20'b00110000110101001010: color_data = 12'b111011101110;
20'b00110000110101001011: color_data = 12'b111011101110;
20'b00110000110101001100: color_data = 12'b111011101110;
20'b00110000110101001101: color_data = 12'b111011101110;
20'b00110000110101001110: color_data = 12'b111011101110;
20'b00110000110101001111: color_data = 12'b111011101110;
20'b00110000110101010001: color_data = 12'b111011101110;
20'b00110000110101010010: color_data = 12'b111011101110;
20'b00110000110101010011: color_data = 12'b111011101110;
20'b00110000110101010100: color_data = 12'b111011101110;
20'b00110000110101010101: color_data = 12'b111011101110;
20'b00110000110101010110: color_data = 12'b111011101110;
20'b00110000110101010111: color_data = 12'b111011101110;
20'b00110000110101011000: color_data = 12'b111011101110;
20'b00110000110101011001: color_data = 12'b111011101110;
20'b00110000110101011010: color_data = 12'b111011101110;
20'b00110000110101111101: color_data = 12'b111011101110;
20'b00110000110101111110: color_data = 12'b111011101110;
20'b00110000110101111111: color_data = 12'b111011101110;
20'b00110000110110000000: color_data = 12'b111011101110;
20'b00110000110110000001: color_data = 12'b111011101110;
20'b00110000110110000010: color_data = 12'b111011101110;
20'b00110000110110000011: color_data = 12'b111011101110;
20'b00110000110110000100: color_data = 12'b111011101110;
20'b00110000110110000101: color_data = 12'b111011101110;
20'b00110000110110000110: color_data = 12'b111011101110;
20'b00110000110110001000: color_data = 12'b111011101110;
20'b00110000110110001001: color_data = 12'b111011101110;
20'b00110000110110001010: color_data = 12'b111011101110;
20'b00110000110110001011: color_data = 12'b111011101110;
20'b00110000110110001100: color_data = 12'b111011101110;
20'b00110000110110001101: color_data = 12'b111011101110;
20'b00110000110110001110: color_data = 12'b111011101110;
20'b00110000110110001111: color_data = 12'b111011101110;
20'b00110000110110010000: color_data = 12'b111011101110;
20'b00110000110110010001: color_data = 12'b111011101110;
20'b00110000110110011110: color_data = 12'b111011101110;
20'b00110000110110011111: color_data = 12'b111011101110;
20'b00110000110110100000: color_data = 12'b111011101110;
20'b00110000110110100001: color_data = 12'b111011101110;
20'b00110000110110100010: color_data = 12'b111011101110;
20'b00110000110110100011: color_data = 12'b111011101110;
20'b00110000110110100100: color_data = 12'b111011101110;
20'b00110000110110100101: color_data = 12'b111011101110;
20'b00110000110110100110: color_data = 12'b111011101110;
20'b00110000110110100111: color_data = 12'b111011101110;
20'b00110000110110101001: color_data = 12'b111011101110;
20'b00110000110110101010: color_data = 12'b111011101110;
20'b00110000110110101011: color_data = 12'b111011101110;
20'b00110000110110101100: color_data = 12'b111011101110;
20'b00110000110110101101: color_data = 12'b111011101110;
20'b00110000110110101110: color_data = 12'b111011101110;
20'b00110000110110101111: color_data = 12'b111011101110;
20'b00110000110110110000: color_data = 12'b111011101110;
20'b00110000110110110001: color_data = 12'b111011101110;
20'b00110000110110110010: color_data = 12'b111011101110;
20'b00110000110110110100: color_data = 12'b111011101110;
20'b00110000110110110101: color_data = 12'b111011101110;
20'b00110000110110110110: color_data = 12'b111011101110;
20'b00110000110110110111: color_data = 12'b111011101110;
20'b00110000110110111000: color_data = 12'b111011101110;
20'b00110000110110111001: color_data = 12'b111011101110;
20'b00110000110110111010: color_data = 12'b111011101110;
20'b00110000110110111011: color_data = 12'b111011101110;
20'b00110000110110111100: color_data = 12'b111011101110;
20'b00110000110110111101: color_data = 12'b111011101110;
20'b00110000110110111111: color_data = 12'b111011101110;
20'b00110000110111000000: color_data = 12'b111011101110;
20'b00110000110111000001: color_data = 12'b111011101110;
20'b00110000110111000010: color_data = 12'b111011101110;
20'b00110000110111000011: color_data = 12'b111011101110;
20'b00110000110111000100: color_data = 12'b111011101110;
20'b00110000110111000101: color_data = 12'b111011101110;
20'b00110000110111000110: color_data = 12'b111011101110;
20'b00110000110111000111: color_data = 12'b111011101110;
20'b00110000110111001000: color_data = 12'b111011101110;
20'b00110000110111001010: color_data = 12'b111011101110;
20'b00110000110111001011: color_data = 12'b111011101110;
20'b00110000110111001100: color_data = 12'b111011101110;
20'b00110000110111001101: color_data = 12'b111011101110;
20'b00110000110111001110: color_data = 12'b111011101110;
20'b00110000110111001111: color_data = 12'b111011101110;
20'b00110000110111010000: color_data = 12'b111011101110;
20'b00110000110111010001: color_data = 12'b111011101110;
20'b00110000110111010010: color_data = 12'b111011101110;
20'b00110000110111010011: color_data = 12'b111011101110;
20'b00110000110111010101: color_data = 12'b111011101110;
20'b00110000110111010110: color_data = 12'b111011101110;
20'b00110000110111010111: color_data = 12'b111011101110;
20'b00110000110111011000: color_data = 12'b111011101110;
20'b00110000110111011001: color_data = 12'b111011101110;
20'b00110000110111011010: color_data = 12'b111011101110;
20'b00110000110111011011: color_data = 12'b111011101110;
20'b00110000110111011100: color_data = 12'b111011101110;
20'b00110000110111011101: color_data = 12'b111011101110;
20'b00110000110111011110: color_data = 12'b111011101110;
20'b00110000110111100000: color_data = 12'b111011101110;
20'b00110000110111100001: color_data = 12'b111011101110;
20'b00110000110111100010: color_data = 12'b111011101110;
20'b00110000110111100011: color_data = 12'b111011101110;
20'b00110000110111100100: color_data = 12'b111011101110;
20'b00110000110111100101: color_data = 12'b111011101110;
20'b00110000110111100110: color_data = 12'b111011101110;
20'b00110000110111100111: color_data = 12'b111011101110;
20'b00110000110111101000: color_data = 12'b111011101110;
20'b00110000110111101001: color_data = 12'b111011101110;
20'b00110001000010100001: color_data = 12'b111011101110;
20'b00110001000010100010: color_data = 12'b111011101110;
20'b00110001000010100011: color_data = 12'b111011101110;
20'b00110001000010100100: color_data = 12'b111011101110;
20'b00110001000010100101: color_data = 12'b111011101110;
20'b00110001000010100110: color_data = 12'b111011101110;
20'b00110001000010100111: color_data = 12'b111011101110;
20'b00110001000010101000: color_data = 12'b111011101110;
20'b00110001000010101001: color_data = 12'b111011101110;
20'b00110001000010101010: color_data = 12'b111011101110;
20'b00110001000010101100: color_data = 12'b111011101110;
20'b00110001000010101101: color_data = 12'b111011101110;
20'b00110001000010101110: color_data = 12'b111011101110;
20'b00110001000010101111: color_data = 12'b111011101110;
20'b00110001000010110000: color_data = 12'b111011101110;
20'b00110001000010110001: color_data = 12'b111011101110;
20'b00110001000010110010: color_data = 12'b111011101110;
20'b00110001000010110011: color_data = 12'b111011101110;
20'b00110001000010110100: color_data = 12'b111011101110;
20'b00110001000010110101: color_data = 12'b111011101110;
20'b00110001000010110111: color_data = 12'b111011101110;
20'b00110001000010111000: color_data = 12'b111011101110;
20'b00110001000010111001: color_data = 12'b111011101110;
20'b00110001000010111010: color_data = 12'b111011101110;
20'b00110001000010111011: color_data = 12'b111011101110;
20'b00110001000010111100: color_data = 12'b111011101110;
20'b00110001000010111101: color_data = 12'b111011101110;
20'b00110001000010111110: color_data = 12'b111011101110;
20'b00110001000010111111: color_data = 12'b111011101110;
20'b00110001000011000000: color_data = 12'b111011101110;
20'b00110001000011000010: color_data = 12'b111011101110;
20'b00110001000011000011: color_data = 12'b111011101110;
20'b00110001000011000100: color_data = 12'b111011101110;
20'b00110001000011000101: color_data = 12'b111011101110;
20'b00110001000011000110: color_data = 12'b111011101110;
20'b00110001000011000111: color_data = 12'b111011101110;
20'b00110001000011001000: color_data = 12'b111011101110;
20'b00110001000011001001: color_data = 12'b111011101110;
20'b00110001000011001010: color_data = 12'b111011101110;
20'b00110001000011001011: color_data = 12'b111011101110;
20'b00110001000011001101: color_data = 12'b111011101110;
20'b00110001000011001110: color_data = 12'b111011101110;
20'b00110001000011001111: color_data = 12'b111011101110;
20'b00110001000011010000: color_data = 12'b111011101110;
20'b00110001000011010001: color_data = 12'b111011101110;
20'b00110001000011010010: color_data = 12'b111011101110;
20'b00110001000011010011: color_data = 12'b111011101110;
20'b00110001000011010100: color_data = 12'b111011101110;
20'b00110001000011010101: color_data = 12'b111011101110;
20'b00110001000011010110: color_data = 12'b111011101110;
20'b00110001000011101110: color_data = 12'b111011101110;
20'b00110001000011101111: color_data = 12'b111011101110;
20'b00110001000011110000: color_data = 12'b111011101110;
20'b00110001000011110001: color_data = 12'b111011101110;
20'b00110001000011110010: color_data = 12'b111011101110;
20'b00110001000011110011: color_data = 12'b111011101110;
20'b00110001000011110100: color_data = 12'b111011101110;
20'b00110001000011110101: color_data = 12'b111011101110;
20'b00110001000011110110: color_data = 12'b111011101110;
20'b00110001000011110111: color_data = 12'b111011101110;
20'b00110001000011111001: color_data = 12'b111011101110;
20'b00110001000011111010: color_data = 12'b111011101110;
20'b00110001000011111011: color_data = 12'b111011101110;
20'b00110001000011111100: color_data = 12'b111011101110;
20'b00110001000011111101: color_data = 12'b111011101110;
20'b00110001000011111110: color_data = 12'b111011101110;
20'b00110001000011111111: color_data = 12'b111011101110;
20'b00110001000100000000: color_data = 12'b111011101110;
20'b00110001000100000001: color_data = 12'b111011101110;
20'b00110001000100000010: color_data = 12'b111011101110;
20'b00110001000100100101: color_data = 12'b111011101110;
20'b00110001000100100110: color_data = 12'b111011101110;
20'b00110001000100100111: color_data = 12'b111011101110;
20'b00110001000100101000: color_data = 12'b111011101110;
20'b00110001000100101001: color_data = 12'b111011101110;
20'b00110001000100101010: color_data = 12'b111011101110;
20'b00110001000100101011: color_data = 12'b111011101110;
20'b00110001000100101100: color_data = 12'b111011101110;
20'b00110001000100101101: color_data = 12'b111011101110;
20'b00110001000100101110: color_data = 12'b111011101110;
20'b00110001000100110000: color_data = 12'b111011101110;
20'b00110001000100110001: color_data = 12'b111011101110;
20'b00110001000100110010: color_data = 12'b111011101110;
20'b00110001000100110011: color_data = 12'b111011101110;
20'b00110001000100110100: color_data = 12'b111011101110;
20'b00110001000100110101: color_data = 12'b111011101110;
20'b00110001000100110110: color_data = 12'b111011101110;
20'b00110001000100110111: color_data = 12'b111011101110;
20'b00110001000100111000: color_data = 12'b111011101110;
20'b00110001000100111001: color_data = 12'b111011101110;
20'b00110001000101000110: color_data = 12'b111011101110;
20'b00110001000101000111: color_data = 12'b111011101110;
20'b00110001000101001000: color_data = 12'b111011101110;
20'b00110001000101001001: color_data = 12'b111011101110;
20'b00110001000101001010: color_data = 12'b111011101110;
20'b00110001000101001011: color_data = 12'b111011101110;
20'b00110001000101001100: color_data = 12'b111011101110;
20'b00110001000101001101: color_data = 12'b111011101110;
20'b00110001000101001110: color_data = 12'b111011101110;
20'b00110001000101001111: color_data = 12'b111011101110;
20'b00110001000101010001: color_data = 12'b111011101110;
20'b00110001000101010010: color_data = 12'b111011101110;
20'b00110001000101010011: color_data = 12'b111011101110;
20'b00110001000101010100: color_data = 12'b111011101110;
20'b00110001000101010101: color_data = 12'b111011101110;
20'b00110001000101010110: color_data = 12'b111011101110;
20'b00110001000101010111: color_data = 12'b111011101110;
20'b00110001000101011000: color_data = 12'b111011101110;
20'b00110001000101011001: color_data = 12'b111011101110;
20'b00110001000101011010: color_data = 12'b111011101110;
20'b00110001000101111101: color_data = 12'b111011101110;
20'b00110001000101111110: color_data = 12'b111011101110;
20'b00110001000101111111: color_data = 12'b111011101110;
20'b00110001000110000000: color_data = 12'b111011101110;
20'b00110001000110000001: color_data = 12'b111011101110;
20'b00110001000110000010: color_data = 12'b111011101110;
20'b00110001000110000011: color_data = 12'b111011101110;
20'b00110001000110000100: color_data = 12'b111011101110;
20'b00110001000110000101: color_data = 12'b111011101110;
20'b00110001000110000110: color_data = 12'b111011101110;
20'b00110001000110001000: color_data = 12'b111011101110;
20'b00110001000110001001: color_data = 12'b111011101110;
20'b00110001000110001010: color_data = 12'b111011101110;
20'b00110001000110001011: color_data = 12'b111011101110;
20'b00110001000110001100: color_data = 12'b111011101110;
20'b00110001000110001101: color_data = 12'b111011101110;
20'b00110001000110001110: color_data = 12'b111011101110;
20'b00110001000110001111: color_data = 12'b111011101110;
20'b00110001000110010000: color_data = 12'b111011101110;
20'b00110001000110010001: color_data = 12'b111011101110;
20'b00110001000110011110: color_data = 12'b111011101110;
20'b00110001000110011111: color_data = 12'b111011101110;
20'b00110001000110100000: color_data = 12'b111011101110;
20'b00110001000110100001: color_data = 12'b111011101110;
20'b00110001000110100010: color_data = 12'b111011101110;
20'b00110001000110100011: color_data = 12'b111011101110;
20'b00110001000110100100: color_data = 12'b111011101110;
20'b00110001000110100101: color_data = 12'b111011101110;
20'b00110001000110100110: color_data = 12'b111011101110;
20'b00110001000110100111: color_data = 12'b111011101110;
20'b00110001000110101001: color_data = 12'b111011101110;
20'b00110001000110101010: color_data = 12'b111011101110;
20'b00110001000110101011: color_data = 12'b111011101110;
20'b00110001000110101100: color_data = 12'b111011101110;
20'b00110001000110101101: color_data = 12'b111011101110;
20'b00110001000110101110: color_data = 12'b111011101110;
20'b00110001000110101111: color_data = 12'b111011101110;
20'b00110001000110110000: color_data = 12'b111011101110;
20'b00110001000110110001: color_data = 12'b111011101110;
20'b00110001000110110010: color_data = 12'b111011101110;
20'b00110001000110110100: color_data = 12'b111011101110;
20'b00110001000110110101: color_data = 12'b111011101110;
20'b00110001000110110110: color_data = 12'b111011101110;
20'b00110001000110110111: color_data = 12'b111011101110;
20'b00110001000110111000: color_data = 12'b111011101110;
20'b00110001000110111001: color_data = 12'b111011101110;
20'b00110001000110111010: color_data = 12'b111011101110;
20'b00110001000110111011: color_data = 12'b111011101110;
20'b00110001000110111100: color_data = 12'b111011101110;
20'b00110001000110111101: color_data = 12'b111011101110;
20'b00110001000110111111: color_data = 12'b111011101110;
20'b00110001000111000000: color_data = 12'b111011101110;
20'b00110001000111000001: color_data = 12'b111011101110;
20'b00110001000111000010: color_data = 12'b111011101110;
20'b00110001000111000011: color_data = 12'b111011101110;
20'b00110001000111000100: color_data = 12'b111011101110;
20'b00110001000111000101: color_data = 12'b111011101110;
20'b00110001000111000110: color_data = 12'b111011101110;
20'b00110001000111000111: color_data = 12'b111011101110;
20'b00110001000111001000: color_data = 12'b111011101110;
20'b00110001000111001010: color_data = 12'b111011101110;
20'b00110001000111001011: color_data = 12'b111011101110;
20'b00110001000111001100: color_data = 12'b111011101110;
20'b00110001000111001101: color_data = 12'b111011101110;
20'b00110001000111001110: color_data = 12'b111011101110;
20'b00110001000111001111: color_data = 12'b111011101110;
20'b00110001000111010000: color_data = 12'b111011101110;
20'b00110001000111010001: color_data = 12'b111011101110;
20'b00110001000111010010: color_data = 12'b111011101110;
20'b00110001000111010011: color_data = 12'b111011101110;
20'b00110001000111010101: color_data = 12'b111011101110;
20'b00110001000111010110: color_data = 12'b111011101110;
20'b00110001000111010111: color_data = 12'b111011101110;
20'b00110001000111011000: color_data = 12'b111011101110;
20'b00110001000111011001: color_data = 12'b111011101110;
20'b00110001000111011010: color_data = 12'b111011101110;
20'b00110001000111011011: color_data = 12'b111011101110;
20'b00110001000111011100: color_data = 12'b111011101110;
20'b00110001000111011101: color_data = 12'b111011101110;
20'b00110001000111011110: color_data = 12'b111011101110;
20'b00110001000111100000: color_data = 12'b111011101110;
20'b00110001000111100001: color_data = 12'b111011101110;
20'b00110001000111100010: color_data = 12'b111011101110;
20'b00110001000111100011: color_data = 12'b111011101110;
20'b00110001000111100100: color_data = 12'b111011101110;
20'b00110001000111100101: color_data = 12'b111011101110;
20'b00110001000111100110: color_data = 12'b111011101110;
20'b00110001000111100111: color_data = 12'b111011101110;
20'b00110001000111101000: color_data = 12'b111011101110;
20'b00110001000111101001: color_data = 12'b111011101110;
20'b00110001010010100001: color_data = 12'b111011101110;
20'b00110001010010100010: color_data = 12'b111011101110;
20'b00110001010010100011: color_data = 12'b111011101110;
20'b00110001010010100100: color_data = 12'b111011101110;
20'b00110001010010100101: color_data = 12'b111011101110;
20'b00110001010010100110: color_data = 12'b111011101110;
20'b00110001010010100111: color_data = 12'b111011101110;
20'b00110001010010101000: color_data = 12'b111011101110;
20'b00110001010010101001: color_data = 12'b111011101110;
20'b00110001010010101010: color_data = 12'b111011101110;
20'b00110001010010101100: color_data = 12'b111011101110;
20'b00110001010010101101: color_data = 12'b111011101110;
20'b00110001010010101110: color_data = 12'b111011101110;
20'b00110001010010101111: color_data = 12'b111011101110;
20'b00110001010010110000: color_data = 12'b111011101110;
20'b00110001010010110001: color_data = 12'b111011101110;
20'b00110001010010110010: color_data = 12'b111011101110;
20'b00110001010010110011: color_data = 12'b111011101110;
20'b00110001010010110100: color_data = 12'b111011101110;
20'b00110001010010110101: color_data = 12'b111011101110;
20'b00110001010010110111: color_data = 12'b111011101110;
20'b00110001010010111000: color_data = 12'b111011101110;
20'b00110001010010111001: color_data = 12'b111011101110;
20'b00110001010010111010: color_data = 12'b111011101110;
20'b00110001010010111011: color_data = 12'b111011101110;
20'b00110001010010111100: color_data = 12'b111011101110;
20'b00110001010010111101: color_data = 12'b111011101110;
20'b00110001010010111110: color_data = 12'b111011101110;
20'b00110001010010111111: color_data = 12'b111011101110;
20'b00110001010011000000: color_data = 12'b111011101110;
20'b00110001010011000010: color_data = 12'b111011101110;
20'b00110001010011000011: color_data = 12'b111011101110;
20'b00110001010011000100: color_data = 12'b111011101110;
20'b00110001010011000101: color_data = 12'b111011101110;
20'b00110001010011000110: color_data = 12'b111011101110;
20'b00110001010011000111: color_data = 12'b111011101110;
20'b00110001010011001000: color_data = 12'b111011101110;
20'b00110001010011001001: color_data = 12'b111011101110;
20'b00110001010011001010: color_data = 12'b111011101110;
20'b00110001010011001011: color_data = 12'b111011101110;
20'b00110001010011001101: color_data = 12'b111011101110;
20'b00110001010011001110: color_data = 12'b111011101110;
20'b00110001010011001111: color_data = 12'b111011101110;
20'b00110001010011010000: color_data = 12'b111011101110;
20'b00110001010011010001: color_data = 12'b111011101110;
20'b00110001010011010010: color_data = 12'b111011101110;
20'b00110001010011010011: color_data = 12'b111011101110;
20'b00110001010011010100: color_data = 12'b111011101110;
20'b00110001010011010101: color_data = 12'b111011101110;
20'b00110001010011010110: color_data = 12'b111011101110;
20'b00110001010011101110: color_data = 12'b111011101110;
20'b00110001010011101111: color_data = 12'b111011101110;
20'b00110001010011110000: color_data = 12'b111011101110;
20'b00110001010011110001: color_data = 12'b111011101110;
20'b00110001010011110010: color_data = 12'b111011101110;
20'b00110001010011110011: color_data = 12'b111011101110;
20'b00110001010011110100: color_data = 12'b111011101110;
20'b00110001010011110101: color_data = 12'b111011101110;
20'b00110001010011110110: color_data = 12'b111011101110;
20'b00110001010011110111: color_data = 12'b111011101110;
20'b00110001010011111001: color_data = 12'b111011101110;
20'b00110001010011111010: color_data = 12'b111011101110;
20'b00110001010011111011: color_data = 12'b111011101110;
20'b00110001010011111100: color_data = 12'b111011101110;
20'b00110001010011111101: color_data = 12'b111011101110;
20'b00110001010011111110: color_data = 12'b111011101110;
20'b00110001010011111111: color_data = 12'b111011101110;
20'b00110001010100000000: color_data = 12'b111011101110;
20'b00110001010100000001: color_data = 12'b111011101110;
20'b00110001010100000010: color_data = 12'b111011101110;
20'b00110001010100100101: color_data = 12'b111011101110;
20'b00110001010100100110: color_data = 12'b111011101110;
20'b00110001010100100111: color_data = 12'b111011101110;
20'b00110001010100101000: color_data = 12'b111011101110;
20'b00110001010100101001: color_data = 12'b111011101110;
20'b00110001010100101010: color_data = 12'b111011101110;
20'b00110001010100101011: color_data = 12'b111011101110;
20'b00110001010100101100: color_data = 12'b111011101110;
20'b00110001010100101101: color_data = 12'b111011101110;
20'b00110001010100101110: color_data = 12'b111011101110;
20'b00110001010100110000: color_data = 12'b111011101110;
20'b00110001010100110001: color_data = 12'b111011101110;
20'b00110001010100110010: color_data = 12'b111011101110;
20'b00110001010100110011: color_data = 12'b111011101110;
20'b00110001010100110100: color_data = 12'b111011101110;
20'b00110001010100110101: color_data = 12'b111011101110;
20'b00110001010100110110: color_data = 12'b111011101110;
20'b00110001010100110111: color_data = 12'b111011101110;
20'b00110001010100111000: color_data = 12'b111011101110;
20'b00110001010100111001: color_data = 12'b111011101110;
20'b00110001010101000110: color_data = 12'b111011101110;
20'b00110001010101000111: color_data = 12'b111011101110;
20'b00110001010101001000: color_data = 12'b111011101110;
20'b00110001010101001001: color_data = 12'b111011101110;
20'b00110001010101001010: color_data = 12'b111011101110;
20'b00110001010101001011: color_data = 12'b111011101110;
20'b00110001010101001100: color_data = 12'b111011101110;
20'b00110001010101001101: color_data = 12'b111011101110;
20'b00110001010101001110: color_data = 12'b111011101110;
20'b00110001010101001111: color_data = 12'b111011101110;
20'b00110001010101010001: color_data = 12'b111011101110;
20'b00110001010101010010: color_data = 12'b111011101110;
20'b00110001010101010011: color_data = 12'b111011101110;
20'b00110001010101010100: color_data = 12'b111011101110;
20'b00110001010101010101: color_data = 12'b111011101110;
20'b00110001010101010110: color_data = 12'b111011101110;
20'b00110001010101010111: color_data = 12'b111011101110;
20'b00110001010101011000: color_data = 12'b111011101110;
20'b00110001010101011001: color_data = 12'b111011101110;
20'b00110001010101011010: color_data = 12'b111011101110;
20'b00110001010101111101: color_data = 12'b111011101110;
20'b00110001010101111110: color_data = 12'b111011101110;
20'b00110001010101111111: color_data = 12'b111011101110;
20'b00110001010110000000: color_data = 12'b111011101110;
20'b00110001010110000001: color_data = 12'b111011101110;
20'b00110001010110000010: color_data = 12'b111011101110;
20'b00110001010110000011: color_data = 12'b111011101110;
20'b00110001010110000100: color_data = 12'b111011101110;
20'b00110001010110000101: color_data = 12'b111011101110;
20'b00110001010110000110: color_data = 12'b111011101110;
20'b00110001010110001000: color_data = 12'b111011101110;
20'b00110001010110001001: color_data = 12'b111011101110;
20'b00110001010110001010: color_data = 12'b111011101110;
20'b00110001010110001011: color_data = 12'b111011101110;
20'b00110001010110001100: color_data = 12'b111011101110;
20'b00110001010110001101: color_data = 12'b111011101110;
20'b00110001010110001110: color_data = 12'b111011101110;
20'b00110001010110001111: color_data = 12'b111011101110;
20'b00110001010110010000: color_data = 12'b111011101110;
20'b00110001010110010001: color_data = 12'b111011101110;
20'b00110001010110011110: color_data = 12'b111011101110;
20'b00110001010110011111: color_data = 12'b111011101110;
20'b00110001010110100000: color_data = 12'b111011101110;
20'b00110001010110100001: color_data = 12'b111011101110;
20'b00110001010110100010: color_data = 12'b111011101110;
20'b00110001010110100011: color_data = 12'b111011101110;
20'b00110001010110100100: color_data = 12'b111011101110;
20'b00110001010110100101: color_data = 12'b111011101110;
20'b00110001010110100110: color_data = 12'b111011101110;
20'b00110001010110100111: color_data = 12'b111011101110;
20'b00110001010110101001: color_data = 12'b111011101110;
20'b00110001010110101010: color_data = 12'b111011101110;
20'b00110001010110101011: color_data = 12'b111011101110;
20'b00110001010110101100: color_data = 12'b111011101110;
20'b00110001010110101101: color_data = 12'b111011101110;
20'b00110001010110101110: color_data = 12'b111011101110;
20'b00110001010110101111: color_data = 12'b111011101110;
20'b00110001010110110000: color_data = 12'b111011101110;
20'b00110001010110110001: color_data = 12'b111011101110;
20'b00110001010110110010: color_data = 12'b111011101110;
20'b00110001010110110100: color_data = 12'b111011101110;
20'b00110001010110110101: color_data = 12'b111011101110;
20'b00110001010110110110: color_data = 12'b111011101110;
20'b00110001010110110111: color_data = 12'b111011101110;
20'b00110001010110111000: color_data = 12'b111011101110;
20'b00110001010110111001: color_data = 12'b111011101110;
20'b00110001010110111010: color_data = 12'b111011101110;
20'b00110001010110111011: color_data = 12'b111011101110;
20'b00110001010110111100: color_data = 12'b111011101110;
20'b00110001010110111101: color_data = 12'b111011101110;
20'b00110001010110111111: color_data = 12'b111011101110;
20'b00110001010111000000: color_data = 12'b111011101110;
20'b00110001010111000001: color_data = 12'b111011101110;
20'b00110001010111000010: color_data = 12'b111011101110;
20'b00110001010111000011: color_data = 12'b111011101110;
20'b00110001010111000100: color_data = 12'b111011101110;
20'b00110001010111000101: color_data = 12'b111011101110;
20'b00110001010111000110: color_data = 12'b111011101110;
20'b00110001010111000111: color_data = 12'b111011101110;
20'b00110001010111001000: color_data = 12'b111011101110;
20'b00110001010111001010: color_data = 12'b111011101110;
20'b00110001010111001011: color_data = 12'b111011101110;
20'b00110001010111001100: color_data = 12'b111011101110;
20'b00110001010111001101: color_data = 12'b111011101110;
20'b00110001010111001110: color_data = 12'b111011101110;
20'b00110001010111001111: color_data = 12'b111011101110;
20'b00110001010111010000: color_data = 12'b111011101110;
20'b00110001010111010001: color_data = 12'b111011101110;
20'b00110001010111010010: color_data = 12'b111011101110;
20'b00110001010111010011: color_data = 12'b111011101110;
20'b00110001010111010101: color_data = 12'b111011101110;
20'b00110001010111010110: color_data = 12'b111011101110;
20'b00110001010111010111: color_data = 12'b111011101110;
20'b00110001010111011000: color_data = 12'b111011101110;
20'b00110001010111011001: color_data = 12'b111011101110;
20'b00110001010111011010: color_data = 12'b111011101110;
20'b00110001010111011011: color_data = 12'b111011101110;
20'b00110001010111011100: color_data = 12'b111011101110;
20'b00110001010111011101: color_data = 12'b111011101110;
20'b00110001010111011110: color_data = 12'b111011101110;
20'b00110001010111100000: color_data = 12'b111011101110;
20'b00110001010111100001: color_data = 12'b111011101110;
20'b00110001010111100010: color_data = 12'b111011101110;
20'b00110001010111100011: color_data = 12'b111011101110;
20'b00110001010111100100: color_data = 12'b111011101110;
20'b00110001010111100101: color_data = 12'b111011101110;
20'b00110001010111100110: color_data = 12'b111011101110;
20'b00110001010111100111: color_data = 12'b111011101110;
20'b00110001010111101000: color_data = 12'b111011101110;
20'b00110001010111101001: color_data = 12'b111011101110;
20'b00111010100010100001: color_data = 12'b111100001111;
20'b00111010100010100010: color_data = 12'b111100001111;
20'b00111010100010100011: color_data = 12'b111100001111;
20'b00111010100010100100: color_data = 12'b111100001111;
20'b00111010100010100101: color_data = 12'b111100001111;
20'b00111010100010100110: color_data = 12'b111100001111;
20'b00111010100010100111: color_data = 12'b111100001111;
20'b00111010100010101000: color_data = 12'b111100001111;
20'b00111010100010101001: color_data = 12'b111100001111;
20'b00111010100010101010: color_data = 12'b111100001111;
20'b00111010100010101100: color_data = 12'b111100001111;
20'b00111010100010101101: color_data = 12'b111100001111;
20'b00111010100010101110: color_data = 12'b111100001111;
20'b00111010100010101111: color_data = 12'b111100001111;
20'b00111010100010110000: color_data = 12'b111100001111;
20'b00111010100010110001: color_data = 12'b111100001111;
20'b00111010100010110010: color_data = 12'b111100001111;
20'b00111010100010110011: color_data = 12'b111100001111;
20'b00111010100010110100: color_data = 12'b111100001111;
20'b00111010100010110101: color_data = 12'b111100001111;
20'b00111010100100100100: color_data = 12'b001111111111;
20'b00111010100100100101: color_data = 12'b001111111111;
20'b00111010100100100110: color_data = 12'b001111111111;
20'b00111010100100100111: color_data = 12'b001111111111;
20'b00111010100100101000: color_data = 12'b001111111111;
20'b00111010100100101001: color_data = 12'b001111111111;
20'b00111010100100101010: color_data = 12'b001111111111;
20'b00111010100100101011: color_data = 12'b001111111111;
20'b00111010100100101100: color_data = 12'b001111111111;
20'b00111010100100101101: color_data = 12'b001111111111;
20'b00111010100100101111: color_data = 12'b001111111111;
20'b00111010100100110000: color_data = 12'b001111111111;
20'b00111010100100110001: color_data = 12'b001111111111;
20'b00111010100100110010: color_data = 12'b001111111111;
20'b00111010100100110011: color_data = 12'b001111111111;
20'b00111010100100110100: color_data = 12'b001111111111;
20'b00111010100100110101: color_data = 12'b001111111111;
20'b00111010100100110110: color_data = 12'b001111111111;
20'b00111010100100110111: color_data = 12'b001111111111;
20'b00111010100100111000: color_data = 12'b001111111111;
20'b00111010100111010011: color_data = 12'b000000001111;
20'b00111010100111010100: color_data = 12'b000000001111;
20'b00111010100111010101: color_data = 12'b000000001111;
20'b00111010100111010110: color_data = 12'b000000001111;
20'b00111010100111010111: color_data = 12'b000000001111;
20'b00111010100111011000: color_data = 12'b000000001111;
20'b00111010100111011001: color_data = 12'b000000001111;
20'b00111010100111011010: color_data = 12'b000000001111;
20'b00111010100111011011: color_data = 12'b000000001111;
20'b00111010100111011100: color_data = 12'b000000001111;
20'b00111010110010100001: color_data = 12'b111100001111;
20'b00111010110010100010: color_data = 12'b111100001111;
20'b00111010110010100011: color_data = 12'b111100001111;
20'b00111010110010100100: color_data = 12'b111100001111;
20'b00111010110010100101: color_data = 12'b111100001111;
20'b00111010110010100110: color_data = 12'b111100001111;
20'b00111010110010100111: color_data = 12'b111100001111;
20'b00111010110010101000: color_data = 12'b111100001111;
20'b00111010110010101001: color_data = 12'b111100001111;
20'b00111010110010101010: color_data = 12'b111100001111;
20'b00111010110010101100: color_data = 12'b111100001111;
20'b00111010110010101101: color_data = 12'b111100001111;
20'b00111010110010101110: color_data = 12'b111100001111;
20'b00111010110010101111: color_data = 12'b111100001111;
20'b00111010110010110000: color_data = 12'b111100001111;
20'b00111010110010110001: color_data = 12'b111100001111;
20'b00111010110010110010: color_data = 12'b111100001111;
20'b00111010110010110011: color_data = 12'b111100001111;
20'b00111010110010110100: color_data = 12'b111100001111;
20'b00111010110010110101: color_data = 12'b111100001111;
20'b00111010110100100100: color_data = 12'b001111111111;
20'b00111010110100100101: color_data = 12'b001111111111;
20'b00111010110100100110: color_data = 12'b001111111111;
20'b00111010110100100111: color_data = 12'b001111111111;
20'b00111010110100101000: color_data = 12'b001111111111;
20'b00111010110100101001: color_data = 12'b001111111111;
20'b00111010110100101010: color_data = 12'b001111111111;
20'b00111010110100101011: color_data = 12'b001111111111;
20'b00111010110100101100: color_data = 12'b001111111111;
20'b00111010110100101101: color_data = 12'b001111111111;
20'b00111010110100101111: color_data = 12'b001111111111;
20'b00111010110100110000: color_data = 12'b001111111111;
20'b00111010110100110001: color_data = 12'b001111111111;
20'b00111010110100110010: color_data = 12'b001111111111;
20'b00111010110100110011: color_data = 12'b001111111111;
20'b00111010110100110100: color_data = 12'b001111111111;
20'b00111010110100110101: color_data = 12'b001111111111;
20'b00111010110100110110: color_data = 12'b001111111111;
20'b00111010110100110111: color_data = 12'b001111111111;
20'b00111010110100111000: color_data = 12'b001111111111;
20'b00111010110111010011: color_data = 12'b000000001111;
20'b00111010110111010100: color_data = 12'b000000001111;
20'b00111010110111010101: color_data = 12'b000000001111;
20'b00111010110111010110: color_data = 12'b000000001111;
20'b00111010110111010111: color_data = 12'b000000001111;
20'b00111010110111011000: color_data = 12'b000000001111;
20'b00111010110111011001: color_data = 12'b000000001111;
20'b00111010110111011010: color_data = 12'b000000001111;
20'b00111010110111011011: color_data = 12'b000000001111;
20'b00111010110111011100: color_data = 12'b000000001111;
20'b00111011000010100001: color_data = 12'b111100001111;
20'b00111011000010100010: color_data = 12'b111100001111;
20'b00111011000010100011: color_data = 12'b111100001111;
20'b00111011000010100100: color_data = 12'b111100001111;
20'b00111011000010100101: color_data = 12'b111100001111;
20'b00111011000010100110: color_data = 12'b111100001111;
20'b00111011000010100111: color_data = 12'b111100001111;
20'b00111011000010101000: color_data = 12'b111100001111;
20'b00111011000010101001: color_data = 12'b111100001111;
20'b00111011000010101010: color_data = 12'b111100001111;
20'b00111011000010101100: color_data = 12'b111100001111;
20'b00111011000010101101: color_data = 12'b111100001111;
20'b00111011000010101110: color_data = 12'b111100001111;
20'b00111011000010101111: color_data = 12'b111100001111;
20'b00111011000010110000: color_data = 12'b111100001111;
20'b00111011000010110001: color_data = 12'b111100001111;
20'b00111011000010110010: color_data = 12'b111100001111;
20'b00111011000010110011: color_data = 12'b111100001111;
20'b00111011000010110100: color_data = 12'b111100001111;
20'b00111011000010110101: color_data = 12'b111100001111;
20'b00111011000100100100: color_data = 12'b001111111111;
20'b00111011000100100101: color_data = 12'b001111111111;
20'b00111011000100100110: color_data = 12'b001111111111;
20'b00111011000100100111: color_data = 12'b001111111111;
20'b00111011000100101000: color_data = 12'b001111111111;
20'b00111011000100101001: color_data = 12'b001111111111;
20'b00111011000100101010: color_data = 12'b001111111111;
20'b00111011000100101011: color_data = 12'b001111111111;
20'b00111011000100101100: color_data = 12'b001111111111;
20'b00111011000100101101: color_data = 12'b001111111111;
20'b00111011000100101111: color_data = 12'b001111111111;
20'b00111011000100110000: color_data = 12'b001111111111;
20'b00111011000100110001: color_data = 12'b001111111111;
20'b00111011000100110010: color_data = 12'b001111111111;
20'b00111011000100110011: color_data = 12'b001111111111;
20'b00111011000100110100: color_data = 12'b001111111111;
20'b00111011000100110101: color_data = 12'b001111111111;
20'b00111011000100110110: color_data = 12'b001111111111;
20'b00111011000100110111: color_data = 12'b001111111111;
20'b00111011000100111000: color_data = 12'b001111111111;
20'b00111011000111010011: color_data = 12'b000000001111;
20'b00111011000111010100: color_data = 12'b000000001111;
20'b00111011000111010101: color_data = 12'b000000001111;
20'b00111011000111010110: color_data = 12'b000000001111;
20'b00111011000111010111: color_data = 12'b000000001111;
20'b00111011000111011000: color_data = 12'b000000001111;
20'b00111011000111011001: color_data = 12'b000000001111;
20'b00111011000111011010: color_data = 12'b000000001111;
20'b00111011000111011011: color_data = 12'b000000001111;
20'b00111011000111011100: color_data = 12'b000000001111;
20'b00111011010010100001: color_data = 12'b111100001111;
20'b00111011010010100010: color_data = 12'b111100001111;
20'b00111011010010100011: color_data = 12'b111100001111;
20'b00111011010010100100: color_data = 12'b111100001111;
20'b00111011010010100101: color_data = 12'b111100001111;
20'b00111011010010100110: color_data = 12'b111100001111;
20'b00111011010010100111: color_data = 12'b111100001111;
20'b00111011010010101000: color_data = 12'b111100001111;
20'b00111011010010101001: color_data = 12'b111100001111;
20'b00111011010010101010: color_data = 12'b111100001111;
20'b00111011010010101100: color_data = 12'b111100001111;
20'b00111011010010101101: color_data = 12'b111100001111;
20'b00111011010010101110: color_data = 12'b111100001111;
20'b00111011010010101111: color_data = 12'b111100001111;
20'b00111011010010110000: color_data = 12'b111100001111;
20'b00111011010010110001: color_data = 12'b111100001111;
20'b00111011010010110010: color_data = 12'b111100001111;
20'b00111011010010110011: color_data = 12'b111100001111;
20'b00111011010010110100: color_data = 12'b111100001111;
20'b00111011010010110101: color_data = 12'b111100001111;
20'b00111011010100100100: color_data = 12'b001111111111;
20'b00111011010100100101: color_data = 12'b001111111111;
20'b00111011010100100110: color_data = 12'b001111111111;
20'b00111011010100100111: color_data = 12'b001111111111;
20'b00111011010100101000: color_data = 12'b001111111111;
20'b00111011010100101001: color_data = 12'b001111111111;
20'b00111011010100101010: color_data = 12'b001111111111;
20'b00111011010100101011: color_data = 12'b001111111111;
20'b00111011010100101100: color_data = 12'b001111111111;
20'b00111011010100101101: color_data = 12'b001111111111;
20'b00111011010100101111: color_data = 12'b001111111111;
20'b00111011010100110000: color_data = 12'b001111111111;
20'b00111011010100110001: color_data = 12'b001111111111;
20'b00111011010100110010: color_data = 12'b001111111111;
20'b00111011010100110011: color_data = 12'b001111111111;
20'b00111011010100110100: color_data = 12'b001111111111;
20'b00111011010100110101: color_data = 12'b001111111111;
20'b00111011010100110110: color_data = 12'b001111111111;
20'b00111011010100110111: color_data = 12'b001111111111;
20'b00111011010100111000: color_data = 12'b001111111111;
20'b00111011010111010011: color_data = 12'b000000001111;
20'b00111011010111010100: color_data = 12'b000000001111;
20'b00111011010111010101: color_data = 12'b000000001111;
20'b00111011010111010110: color_data = 12'b000000001111;
20'b00111011010111010111: color_data = 12'b000000001111;
20'b00111011010111011000: color_data = 12'b000000001111;
20'b00111011010111011001: color_data = 12'b000000001111;
20'b00111011010111011010: color_data = 12'b000000001111;
20'b00111011010111011011: color_data = 12'b000000001111;
20'b00111011010111011100: color_data = 12'b000000001111;
20'b00111011100010100001: color_data = 12'b111100001111;
20'b00111011100010100010: color_data = 12'b111100001111;
20'b00111011100010100011: color_data = 12'b111100001111;
20'b00111011100010100100: color_data = 12'b111100001111;
20'b00111011100010100101: color_data = 12'b111100001111;
20'b00111011100010100110: color_data = 12'b111100001111;
20'b00111011100010100111: color_data = 12'b111100001111;
20'b00111011100010101000: color_data = 12'b111100001111;
20'b00111011100010101001: color_data = 12'b111100001111;
20'b00111011100010101010: color_data = 12'b111100001111;
20'b00111011100010101100: color_data = 12'b111100001111;
20'b00111011100010101101: color_data = 12'b111100001111;
20'b00111011100010101110: color_data = 12'b111100001111;
20'b00111011100010101111: color_data = 12'b111100001111;
20'b00111011100010110000: color_data = 12'b111100001111;
20'b00111011100010110001: color_data = 12'b111100001111;
20'b00111011100010110010: color_data = 12'b111100001111;
20'b00111011100010110011: color_data = 12'b111100001111;
20'b00111011100010110100: color_data = 12'b111100001111;
20'b00111011100010110101: color_data = 12'b111100001111;
20'b00111011100100100100: color_data = 12'b001111111111;
20'b00111011100100100101: color_data = 12'b001111111111;
20'b00111011100100100110: color_data = 12'b001111111111;
20'b00111011100100100111: color_data = 12'b001111111111;
20'b00111011100100101000: color_data = 12'b001111111111;
20'b00111011100100101001: color_data = 12'b001111111111;
20'b00111011100100101010: color_data = 12'b001111111111;
20'b00111011100100101011: color_data = 12'b001111111111;
20'b00111011100100101100: color_data = 12'b001111111111;
20'b00111011100100101101: color_data = 12'b001111111111;
20'b00111011100100101111: color_data = 12'b001111111111;
20'b00111011100100110000: color_data = 12'b001111111111;
20'b00111011100100110001: color_data = 12'b001111111111;
20'b00111011100100110010: color_data = 12'b001111111111;
20'b00111011100100110011: color_data = 12'b001111111111;
20'b00111011100100110100: color_data = 12'b001111111111;
20'b00111011100100110101: color_data = 12'b001111111111;
20'b00111011100100110110: color_data = 12'b001111111111;
20'b00111011100100110111: color_data = 12'b001111111111;
20'b00111011100100111000: color_data = 12'b001111111111;
20'b00111011100111010011: color_data = 12'b000000001111;
20'b00111011100111010100: color_data = 12'b000000001111;
20'b00111011100111010101: color_data = 12'b000000001111;
20'b00111011100111010110: color_data = 12'b000000001111;
20'b00111011100111010111: color_data = 12'b000000001111;
20'b00111011100111011000: color_data = 12'b000000001111;
20'b00111011100111011001: color_data = 12'b000000001111;
20'b00111011100111011010: color_data = 12'b000000001111;
20'b00111011100111011011: color_data = 12'b000000001111;
20'b00111011100111011100: color_data = 12'b000000001111;
20'b00111011110010100001: color_data = 12'b111100001111;
20'b00111011110010100010: color_data = 12'b111100001111;
20'b00111011110010100011: color_data = 12'b111100001111;
20'b00111011110010100100: color_data = 12'b111100001111;
20'b00111011110010100101: color_data = 12'b111100001111;
20'b00111011110010100110: color_data = 12'b111100001111;
20'b00111011110010100111: color_data = 12'b111100001111;
20'b00111011110010101000: color_data = 12'b111100001111;
20'b00111011110010101001: color_data = 12'b111100001111;
20'b00111011110010101010: color_data = 12'b111100001111;
20'b00111011110010101100: color_data = 12'b111100001111;
20'b00111011110010101101: color_data = 12'b111100001111;
20'b00111011110010101110: color_data = 12'b111100001111;
20'b00111011110010101111: color_data = 12'b111100001111;
20'b00111011110010110000: color_data = 12'b111100001111;
20'b00111011110010110001: color_data = 12'b111100001111;
20'b00111011110010110010: color_data = 12'b111100001111;
20'b00111011110010110011: color_data = 12'b111100001111;
20'b00111011110010110100: color_data = 12'b111100001111;
20'b00111011110010110101: color_data = 12'b111100001111;
20'b00111011110100100100: color_data = 12'b001111111111;
20'b00111011110100100101: color_data = 12'b001111111111;
20'b00111011110100100110: color_data = 12'b001111111111;
20'b00111011110100100111: color_data = 12'b001111111111;
20'b00111011110100101000: color_data = 12'b001111111111;
20'b00111011110100101001: color_data = 12'b001111111111;
20'b00111011110100101010: color_data = 12'b001111111111;
20'b00111011110100101011: color_data = 12'b001111111111;
20'b00111011110100101100: color_data = 12'b001111111111;
20'b00111011110100101101: color_data = 12'b001111111111;
20'b00111011110100101111: color_data = 12'b001111111111;
20'b00111011110100110000: color_data = 12'b001111111111;
20'b00111011110100110001: color_data = 12'b001111111111;
20'b00111011110100110010: color_data = 12'b001111111111;
20'b00111011110100110011: color_data = 12'b001111111111;
20'b00111011110100110100: color_data = 12'b001111111111;
20'b00111011110100110101: color_data = 12'b001111111111;
20'b00111011110100110110: color_data = 12'b001111111111;
20'b00111011110100110111: color_data = 12'b001111111111;
20'b00111011110100111000: color_data = 12'b001111111111;
20'b00111011110111010011: color_data = 12'b000000001111;
20'b00111011110111010100: color_data = 12'b000000001111;
20'b00111011110111010101: color_data = 12'b000000001111;
20'b00111011110111010110: color_data = 12'b000000001111;
20'b00111011110111010111: color_data = 12'b000000001111;
20'b00111011110111011000: color_data = 12'b000000001111;
20'b00111011110111011001: color_data = 12'b000000001111;
20'b00111011110111011010: color_data = 12'b000000001111;
20'b00111011110111011011: color_data = 12'b000000001111;
20'b00111011110111011100: color_data = 12'b000000001111;
20'b00111100000010100001: color_data = 12'b111100001111;
20'b00111100000010100010: color_data = 12'b111100001111;
20'b00111100000010100011: color_data = 12'b111100001111;
20'b00111100000010100100: color_data = 12'b111100001111;
20'b00111100000010100101: color_data = 12'b111100001111;
20'b00111100000010100110: color_data = 12'b111100001111;
20'b00111100000010100111: color_data = 12'b111100001111;
20'b00111100000010101000: color_data = 12'b111100001111;
20'b00111100000010101001: color_data = 12'b111100001111;
20'b00111100000010101010: color_data = 12'b111100001111;
20'b00111100000010101100: color_data = 12'b111100001111;
20'b00111100000010101101: color_data = 12'b111100001111;
20'b00111100000010101110: color_data = 12'b111100001111;
20'b00111100000010101111: color_data = 12'b111100001111;
20'b00111100000010110000: color_data = 12'b111100001111;
20'b00111100000010110001: color_data = 12'b111100001111;
20'b00111100000010110010: color_data = 12'b111100001111;
20'b00111100000010110011: color_data = 12'b111100001111;
20'b00111100000010110100: color_data = 12'b111100001111;
20'b00111100000010110101: color_data = 12'b111100001111;
20'b00111100000100100100: color_data = 12'b001111111111;
20'b00111100000100100101: color_data = 12'b001111111111;
20'b00111100000100100110: color_data = 12'b001111111111;
20'b00111100000100100111: color_data = 12'b001111111111;
20'b00111100000100101000: color_data = 12'b001111111111;
20'b00111100000100101001: color_data = 12'b001111111111;
20'b00111100000100101010: color_data = 12'b001111111111;
20'b00111100000100101011: color_data = 12'b001111111111;
20'b00111100000100101100: color_data = 12'b001111111111;
20'b00111100000100101101: color_data = 12'b001111111111;
20'b00111100000100101111: color_data = 12'b001111111111;
20'b00111100000100110000: color_data = 12'b001111111111;
20'b00111100000100110001: color_data = 12'b001111111111;
20'b00111100000100110010: color_data = 12'b001111111111;
20'b00111100000100110011: color_data = 12'b001111111111;
20'b00111100000100110100: color_data = 12'b001111111111;
20'b00111100000100110101: color_data = 12'b001111111111;
20'b00111100000100110110: color_data = 12'b001111111111;
20'b00111100000100110111: color_data = 12'b001111111111;
20'b00111100000100111000: color_data = 12'b001111111111;
20'b00111100000111010011: color_data = 12'b000000001111;
20'b00111100000111010100: color_data = 12'b000000001111;
20'b00111100000111010101: color_data = 12'b000000001111;
20'b00111100000111010110: color_data = 12'b000000001111;
20'b00111100000111010111: color_data = 12'b000000001111;
20'b00111100000111011000: color_data = 12'b000000001111;
20'b00111100000111011001: color_data = 12'b000000001111;
20'b00111100000111011010: color_data = 12'b000000001111;
20'b00111100000111011011: color_data = 12'b000000001111;
20'b00111100000111011100: color_data = 12'b000000001111;
20'b00111100010010100001: color_data = 12'b111100001111;
20'b00111100010010100010: color_data = 12'b111100001111;
20'b00111100010010100011: color_data = 12'b111100001111;
20'b00111100010010100100: color_data = 12'b111100001111;
20'b00111100010010100101: color_data = 12'b111100001111;
20'b00111100010010100110: color_data = 12'b111100001111;
20'b00111100010010100111: color_data = 12'b111100001111;
20'b00111100010010101000: color_data = 12'b111100001111;
20'b00111100010010101001: color_data = 12'b111100001111;
20'b00111100010010101010: color_data = 12'b111100001111;
20'b00111100010010101100: color_data = 12'b111100001111;
20'b00111100010010101101: color_data = 12'b111100001111;
20'b00111100010010101110: color_data = 12'b111100001111;
20'b00111100010010101111: color_data = 12'b111100001111;
20'b00111100010010110000: color_data = 12'b111100001111;
20'b00111100010010110001: color_data = 12'b111100001111;
20'b00111100010010110010: color_data = 12'b111100001111;
20'b00111100010010110011: color_data = 12'b111100001111;
20'b00111100010010110100: color_data = 12'b111100001111;
20'b00111100010010110101: color_data = 12'b111100001111;
20'b00111100010100100100: color_data = 12'b001111111111;
20'b00111100010100100101: color_data = 12'b001111111111;
20'b00111100010100100110: color_data = 12'b001111111111;
20'b00111100010100100111: color_data = 12'b001111111111;
20'b00111100010100101000: color_data = 12'b001111111111;
20'b00111100010100101001: color_data = 12'b001111111111;
20'b00111100010100101010: color_data = 12'b001111111111;
20'b00111100010100101011: color_data = 12'b001111111111;
20'b00111100010100101100: color_data = 12'b001111111111;
20'b00111100010100101101: color_data = 12'b001111111111;
20'b00111100010100101111: color_data = 12'b001111111111;
20'b00111100010100110000: color_data = 12'b001111111111;
20'b00111100010100110001: color_data = 12'b001111111111;
20'b00111100010100110010: color_data = 12'b001111111111;
20'b00111100010100110011: color_data = 12'b001111111111;
20'b00111100010100110100: color_data = 12'b001111111111;
20'b00111100010100110101: color_data = 12'b001111111111;
20'b00111100010100110110: color_data = 12'b001111111111;
20'b00111100010100110111: color_data = 12'b001111111111;
20'b00111100010100111000: color_data = 12'b001111111111;
20'b00111100010111010011: color_data = 12'b000000001111;
20'b00111100010111010100: color_data = 12'b000000001111;
20'b00111100010111010101: color_data = 12'b000000001111;
20'b00111100010111010110: color_data = 12'b000000001111;
20'b00111100010111010111: color_data = 12'b000000001111;
20'b00111100010111011000: color_data = 12'b000000001111;
20'b00111100010111011001: color_data = 12'b000000001111;
20'b00111100010111011010: color_data = 12'b000000001111;
20'b00111100010111011011: color_data = 12'b000000001111;
20'b00111100010111011100: color_data = 12'b000000001111;
20'b00111100100010100001: color_data = 12'b111100001111;
20'b00111100100010100010: color_data = 12'b111100001111;
20'b00111100100010100011: color_data = 12'b111100001111;
20'b00111100100010100100: color_data = 12'b111100001111;
20'b00111100100010100101: color_data = 12'b111100001111;
20'b00111100100010100110: color_data = 12'b111100001111;
20'b00111100100010100111: color_data = 12'b111100001111;
20'b00111100100010101000: color_data = 12'b111100001111;
20'b00111100100010101001: color_data = 12'b111100001111;
20'b00111100100010101010: color_data = 12'b111100001111;
20'b00111100100010101100: color_data = 12'b111100001111;
20'b00111100100010101101: color_data = 12'b111100001111;
20'b00111100100010101110: color_data = 12'b111100001111;
20'b00111100100010101111: color_data = 12'b111100001111;
20'b00111100100010110000: color_data = 12'b111100001111;
20'b00111100100010110001: color_data = 12'b111100001111;
20'b00111100100010110010: color_data = 12'b111100001111;
20'b00111100100010110011: color_data = 12'b111100001111;
20'b00111100100010110100: color_data = 12'b111100001111;
20'b00111100100010110101: color_data = 12'b111100001111;
20'b00111100100100100100: color_data = 12'b001111111111;
20'b00111100100100100101: color_data = 12'b001111111111;
20'b00111100100100100110: color_data = 12'b001111111111;
20'b00111100100100100111: color_data = 12'b001111111111;
20'b00111100100100101000: color_data = 12'b001111111111;
20'b00111100100100101001: color_data = 12'b001111111111;
20'b00111100100100101010: color_data = 12'b001111111111;
20'b00111100100100101011: color_data = 12'b001111111111;
20'b00111100100100101100: color_data = 12'b001111111111;
20'b00111100100100101101: color_data = 12'b001111111111;
20'b00111100100100101111: color_data = 12'b001111111111;
20'b00111100100100110000: color_data = 12'b001111111111;
20'b00111100100100110001: color_data = 12'b001111111111;
20'b00111100100100110010: color_data = 12'b001111111111;
20'b00111100100100110011: color_data = 12'b001111111111;
20'b00111100100100110100: color_data = 12'b001111111111;
20'b00111100100100110101: color_data = 12'b001111111111;
20'b00111100100100110110: color_data = 12'b001111111111;
20'b00111100100100110111: color_data = 12'b001111111111;
20'b00111100100100111000: color_data = 12'b001111111111;
20'b00111100100111010011: color_data = 12'b000000001111;
20'b00111100100111010100: color_data = 12'b000000001111;
20'b00111100100111010101: color_data = 12'b000000001111;
20'b00111100100111010110: color_data = 12'b000000001111;
20'b00111100100111010111: color_data = 12'b000000001111;
20'b00111100100111011000: color_data = 12'b000000001111;
20'b00111100100111011001: color_data = 12'b000000001111;
20'b00111100100111011010: color_data = 12'b000000001111;
20'b00111100100111011011: color_data = 12'b000000001111;
20'b00111100100111011100: color_data = 12'b000000001111;
20'b00111100110010100001: color_data = 12'b111100001111;
20'b00111100110010100010: color_data = 12'b111100001111;
20'b00111100110010100011: color_data = 12'b111100001111;
20'b00111100110010100100: color_data = 12'b111100001111;
20'b00111100110010100101: color_data = 12'b111100001111;
20'b00111100110010100110: color_data = 12'b111100001111;
20'b00111100110010100111: color_data = 12'b111100001111;
20'b00111100110010101000: color_data = 12'b111100001111;
20'b00111100110010101001: color_data = 12'b111100001111;
20'b00111100110010101010: color_data = 12'b111100001111;
20'b00111100110010101100: color_data = 12'b111100001111;
20'b00111100110010101101: color_data = 12'b111100001111;
20'b00111100110010101110: color_data = 12'b111100001111;
20'b00111100110010101111: color_data = 12'b111100001111;
20'b00111100110010110000: color_data = 12'b111100001111;
20'b00111100110010110001: color_data = 12'b111100001111;
20'b00111100110010110010: color_data = 12'b111100001111;
20'b00111100110010110011: color_data = 12'b111100001111;
20'b00111100110010110100: color_data = 12'b111100001111;
20'b00111100110010110101: color_data = 12'b111100001111;
20'b00111100110100100100: color_data = 12'b001111111111;
20'b00111100110100100101: color_data = 12'b001111111111;
20'b00111100110100100110: color_data = 12'b001111111111;
20'b00111100110100100111: color_data = 12'b001111111111;
20'b00111100110100101000: color_data = 12'b001111111111;
20'b00111100110100101001: color_data = 12'b001111111111;
20'b00111100110100101010: color_data = 12'b001111111111;
20'b00111100110100101011: color_data = 12'b001111111111;
20'b00111100110100101100: color_data = 12'b001111111111;
20'b00111100110100101101: color_data = 12'b001111111111;
20'b00111100110100101111: color_data = 12'b001111111111;
20'b00111100110100110000: color_data = 12'b001111111111;
20'b00111100110100110001: color_data = 12'b001111111111;
20'b00111100110100110010: color_data = 12'b001111111111;
20'b00111100110100110011: color_data = 12'b001111111111;
20'b00111100110100110100: color_data = 12'b001111111111;
20'b00111100110100110101: color_data = 12'b001111111111;
20'b00111100110100110110: color_data = 12'b001111111111;
20'b00111100110100110111: color_data = 12'b001111111111;
20'b00111100110100111000: color_data = 12'b001111111111;
20'b00111100110111010011: color_data = 12'b000000001111;
20'b00111100110111010100: color_data = 12'b000000001111;
20'b00111100110111010101: color_data = 12'b000000001111;
20'b00111100110111010110: color_data = 12'b000000001111;
20'b00111100110111010111: color_data = 12'b000000001111;
20'b00111100110111011000: color_data = 12'b000000001111;
20'b00111100110111011001: color_data = 12'b000000001111;
20'b00111100110111011010: color_data = 12'b000000001111;
20'b00111100110111011011: color_data = 12'b000000001111;
20'b00111100110111011100: color_data = 12'b000000001111;
20'b00111101010010100001: color_data = 12'b111100001111;
20'b00111101010010100010: color_data = 12'b111100001111;
20'b00111101010010100011: color_data = 12'b111100001111;
20'b00111101010010100100: color_data = 12'b111100001111;
20'b00111101010010100101: color_data = 12'b111100001111;
20'b00111101010010100110: color_data = 12'b111100001111;
20'b00111101010010100111: color_data = 12'b111100001111;
20'b00111101010010101000: color_data = 12'b111100001111;
20'b00111101010010101001: color_data = 12'b111100001111;
20'b00111101010010101010: color_data = 12'b111100001111;
20'b00111101010011101101: color_data = 12'b000001111111;
20'b00111101010011101110: color_data = 12'b000001111111;
20'b00111101010011101111: color_data = 12'b000001111111;
20'b00111101010011110000: color_data = 12'b000001111111;
20'b00111101010011110001: color_data = 12'b000001111111;
20'b00111101010011110010: color_data = 12'b000001111111;
20'b00111101010011110011: color_data = 12'b000001111111;
20'b00111101010011110100: color_data = 12'b000001111111;
20'b00111101010011110101: color_data = 12'b000001111111;
20'b00111101010011110110: color_data = 12'b000001111111;
20'b00111101010011111000: color_data = 12'b000001111111;
20'b00111101010011111001: color_data = 12'b000001111111;
20'b00111101010011111010: color_data = 12'b000001111111;
20'b00111101010011111011: color_data = 12'b000001111111;
20'b00111101010011111100: color_data = 12'b000001111111;
20'b00111101010011111101: color_data = 12'b000001111111;
20'b00111101010011111110: color_data = 12'b000001111111;
20'b00111101010011111111: color_data = 12'b000001111111;
20'b00111101010100000000: color_data = 12'b000001111111;
20'b00111101010100000001: color_data = 12'b000001111111;
20'b00111101010100100100: color_data = 12'b001111111111;
20'b00111101010100100101: color_data = 12'b001111111111;
20'b00111101010100100110: color_data = 12'b001111111111;
20'b00111101010100100111: color_data = 12'b001111111111;
20'b00111101010100101000: color_data = 12'b001111111111;
20'b00111101010100101001: color_data = 12'b001111111111;
20'b00111101010100101010: color_data = 12'b001111111111;
20'b00111101010100101011: color_data = 12'b001111111111;
20'b00111101010100101100: color_data = 12'b001111111111;
20'b00111101010100101101: color_data = 12'b001111111111;
20'b00111101010100101111: color_data = 12'b001111111111;
20'b00111101010100110000: color_data = 12'b001111111111;
20'b00111101010100110001: color_data = 12'b001111111111;
20'b00111101010100110010: color_data = 12'b001111111111;
20'b00111101010100110011: color_data = 12'b001111111111;
20'b00111101010100110100: color_data = 12'b001111111111;
20'b00111101010100110101: color_data = 12'b001111111111;
20'b00111101010100110110: color_data = 12'b001111111111;
20'b00111101010100110111: color_data = 12'b001111111111;
20'b00111101010100111000: color_data = 12'b001111111111;
20'b00111101010101000100: color_data = 12'b000011110111;
20'b00111101010101000101: color_data = 12'b000011110111;
20'b00111101010101000110: color_data = 12'b000011110111;
20'b00111101010101000111: color_data = 12'b000011110111;
20'b00111101010101001000: color_data = 12'b000011110111;
20'b00111101010101001001: color_data = 12'b000011110111;
20'b00111101010101001010: color_data = 12'b000011110111;
20'b00111101010101001011: color_data = 12'b000011110111;
20'b00111101010101001100: color_data = 12'b000011110111;
20'b00111101010101001101: color_data = 12'b000011110111;
20'b00111101010101001111: color_data = 12'b000011110111;
20'b00111101010101010000: color_data = 12'b000011110111;
20'b00111101010101010001: color_data = 12'b000011110111;
20'b00111101010101010010: color_data = 12'b000011110111;
20'b00111101010101010011: color_data = 12'b000011110111;
20'b00111101010101010100: color_data = 12'b000011110111;
20'b00111101010101010101: color_data = 12'b000011110111;
20'b00111101010101010110: color_data = 12'b000011110111;
20'b00111101010101010111: color_data = 12'b000011110111;
20'b00111101010101011000: color_data = 12'b000011110111;
20'b00111101010101011010: color_data = 12'b000011110111;
20'b00111101010101011011: color_data = 12'b000011110111;
20'b00111101010101011100: color_data = 12'b000011110111;
20'b00111101010101011101: color_data = 12'b000011110111;
20'b00111101010101011110: color_data = 12'b000011110111;
20'b00111101010101011111: color_data = 12'b000011110111;
20'b00111101010101100000: color_data = 12'b000011110111;
20'b00111101010101100001: color_data = 12'b000011110111;
20'b00111101010101100010: color_data = 12'b000011110111;
20'b00111101010101100011: color_data = 12'b000011110111;
20'b00111101010111010011: color_data = 12'b000000001111;
20'b00111101010111010100: color_data = 12'b000000001111;
20'b00111101010111010101: color_data = 12'b000000001111;
20'b00111101010111010110: color_data = 12'b000000001111;
20'b00111101010111010111: color_data = 12'b000000001111;
20'b00111101010111011000: color_data = 12'b000000001111;
20'b00111101010111011001: color_data = 12'b000000001111;
20'b00111101010111011010: color_data = 12'b000000001111;
20'b00111101010111011011: color_data = 12'b000000001111;
20'b00111101010111011100: color_data = 12'b000000001111;
20'b00111101010111011110: color_data = 12'b000000001111;
20'b00111101010111011111: color_data = 12'b000000001111;
20'b00111101010111100000: color_data = 12'b000000001111;
20'b00111101010111100001: color_data = 12'b000000001111;
20'b00111101010111100010: color_data = 12'b000000001111;
20'b00111101010111100011: color_data = 12'b000000001111;
20'b00111101010111100100: color_data = 12'b000000001111;
20'b00111101010111100101: color_data = 12'b000000001111;
20'b00111101010111100110: color_data = 12'b000000001111;
20'b00111101010111100111: color_data = 12'b000000001111;
20'b00111101100010100001: color_data = 12'b111100001111;
20'b00111101100010100010: color_data = 12'b111100001111;
20'b00111101100010100011: color_data = 12'b111100001111;
20'b00111101100010100100: color_data = 12'b111100001111;
20'b00111101100010100101: color_data = 12'b111100001111;
20'b00111101100010100110: color_data = 12'b111100001111;
20'b00111101100010100111: color_data = 12'b111100001111;
20'b00111101100010101000: color_data = 12'b111100001111;
20'b00111101100010101001: color_data = 12'b111100001111;
20'b00111101100010101010: color_data = 12'b111100001111;
20'b00111101100011101101: color_data = 12'b000001111111;
20'b00111101100011101110: color_data = 12'b000001111111;
20'b00111101100011101111: color_data = 12'b000001111111;
20'b00111101100011110000: color_data = 12'b000001111111;
20'b00111101100011110001: color_data = 12'b000001111111;
20'b00111101100011110010: color_data = 12'b000001111111;
20'b00111101100011110011: color_data = 12'b000001111111;
20'b00111101100011110100: color_data = 12'b000001111111;
20'b00111101100011110101: color_data = 12'b000001111111;
20'b00111101100011110110: color_data = 12'b000001111111;
20'b00111101100011111000: color_data = 12'b000001111111;
20'b00111101100011111001: color_data = 12'b000001111111;
20'b00111101100011111010: color_data = 12'b000001111111;
20'b00111101100011111011: color_data = 12'b000001111111;
20'b00111101100011111100: color_data = 12'b000001111111;
20'b00111101100011111101: color_data = 12'b000001111111;
20'b00111101100011111110: color_data = 12'b000001111111;
20'b00111101100011111111: color_data = 12'b000001111111;
20'b00111101100100000000: color_data = 12'b000001111111;
20'b00111101100100000001: color_data = 12'b000001111111;
20'b00111101100100100100: color_data = 12'b001111111111;
20'b00111101100100100101: color_data = 12'b001111111111;
20'b00111101100100100110: color_data = 12'b001111111111;
20'b00111101100100100111: color_data = 12'b001111111111;
20'b00111101100100101000: color_data = 12'b001111111111;
20'b00111101100100101001: color_data = 12'b001111111111;
20'b00111101100100101010: color_data = 12'b001111111111;
20'b00111101100100101011: color_data = 12'b001111111111;
20'b00111101100100101100: color_data = 12'b001111111111;
20'b00111101100100101101: color_data = 12'b001111111111;
20'b00111101100100101111: color_data = 12'b001111111111;
20'b00111101100100110000: color_data = 12'b001111111111;
20'b00111101100100110001: color_data = 12'b001111111111;
20'b00111101100100110010: color_data = 12'b001111111111;
20'b00111101100100110011: color_data = 12'b001111111111;
20'b00111101100100110100: color_data = 12'b001111111111;
20'b00111101100100110101: color_data = 12'b001111111111;
20'b00111101100100110110: color_data = 12'b001111111111;
20'b00111101100100110111: color_data = 12'b001111111111;
20'b00111101100100111000: color_data = 12'b001111111111;
20'b00111101100101000100: color_data = 12'b000011110111;
20'b00111101100101000101: color_data = 12'b000011110111;
20'b00111101100101000110: color_data = 12'b000011110111;
20'b00111101100101000111: color_data = 12'b000011110111;
20'b00111101100101001000: color_data = 12'b000011110111;
20'b00111101100101001001: color_data = 12'b000011110111;
20'b00111101100101001010: color_data = 12'b000011110111;
20'b00111101100101001011: color_data = 12'b000011110111;
20'b00111101100101001100: color_data = 12'b000011110111;
20'b00111101100101001101: color_data = 12'b000011110111;
20'b00111101100101001111: color_data = 12'b000011110111;
20'b00111101100101010000: color_data = 12'b000011110111;
20'b00111101100101010001: color_data = 12'b000011110111;
20'b00111101100101010010: color_data = 12'b000011110111;
20'b00111101100101010011: color_data = 12'b000011110111;
20'b00111101100101010100: color_data = 12'b000011110111;
20'b00111101100101010101: color_data = 12'b000011110111;
20'b00111101100101010110: color_data = 12'b000011110111;
20'b00111101100101010111: color_data = 12'b000011110111;
20'b00111101100101011000: color_data = 12'b000011110111;
20'b00111101100101011010: color_data = 12'b000011110111;
20'b00111101100101011011: color_data = 12'b000011110111;
20'b00111101100101011100: color_data = 12'b000011110111;
20'b00111101100101011101: color_data = 12'b000011110111;
20'b00111101100101011110: color_data = 12'b000011110111;
20'b00111101100101011111: color_data = 12'b000011110111;
20'b00111101100101100000: color_data = 12'b000011110111;
20'b00111101100101100001: color_data = 12'b000011110111;
20'b00111101100101100010: color_data = 12'b000011110111;
20'b00111101100101100011: color_data = 12'b000011110111;
20'b00111101100111010011: color_data = 12'b000000001111;
20'b00111101100111010100: color_data = 12'b000000001111;
20'b00111101100111010101: color_data = 12'b000000001111;
20'b00111101100111010110: color_data = 12'b000000001111;
20'b00111101100111010111: color_data = 12'b000000001111;
20'b00111101100111011000: color_data = 12'b000000001111;
20'b00111101100111011001: color_data = 12'b000000001111;
20'b00111101100111011010: color_data = 12'b000000001111;
20'b00111101100111011011: color_data = 12'b000000001111;
20'b00111101100111011100: color_data = 12'b000000001111;
20'b00111101100111011110: color_data = 12'b000000001111;
20'b00111101100111011111: color_data = 12'b000000001111;
20'b00111101100111100000: color_data = 12'b000000001111;
20'b00111101100111100001: color_data = 12'b000000001111;
20'b00111101100111100010: color_data = 12'b000000001111;
20'b00111101100111100011: color_data = 12'b000000001111;
20'b00111101100111100100: color_data = 12'b000000001111;
20'b00111101100111100101: color_data = 12'b000000001111;
20'b00111101100111100110: color_data = 12'b000000001111;
20'b00111101100111100111: color_data = 12'b000000001111;
20'b00111101110010100001: color_data = 12'b111100001111;
20'b00111101110010100010: color_data = 12'b111100001111;
20'b00111101110010100011: color_data = 12'b111100001111;
20'b00111101110010100100: color_data = 12'b111100001111;
20'b00111101110010100101: color_data = 12'b111100001111;
20'b00111101110010100110: color_data = 12'b111100001111;
20'b00111101110010100111: color_data = 12'b111100001111;
20'b00111101110010101000: color_data = 12'b111100001111;
20'b00111101110010101001: color_data = 12'b111100001111;
20'b00111101110010101010: color_data = 12'b111100001111;
20'b00111101110011101101: color_data = 12'b000001111111;
20'b00111101110011101110: color_data = 12'b000001111111;
20'b00111101110011101111: color_data = 12'b000001111111;
20'b00111101110011110000: color_data = 12'b000001111111;
20'b00111101110011110001: color_data = 12'b000001111111;
20'b00111101110011110010: color_data = 12'b000001111111;
20'b00111101110011110011: color_data = 12'b000001111111;
20'b00111101110011110100: color_data = 12'b000001111111;
20'b00111101110011110101: color_data = 12'b000001111111;
20'b00111101110011110110: color_data = 12'b000001111111;
20'b00111101110011111000: color_data = 12'b000001111111;
20'b00111101110011111001: color_data = 12'b000001111111;
20'b00111101110011111010: color_data = 12'b000001111111;
20'b00111101110011111011: color_data = 12'b000001111111;
20'b00111101110011111100: color_data = 12'b000001111111;
20'b00111101110011111101: color_data = 12'b000001111111;
20'b00111101110011111110: color_data = 12'b000001111111;
20'b00111101110011111111: color_data = 12'b000001111111;
20'b00111101110100000000: color_data = 12'b000001111111;
20'b00111101110100000001: color_data = 12'b000001111111;
20'b00111101110100100100: color_data = 12'b001111111111;
20'b00111101110100100101: color_data = 12'b001111111111;
20'b00111101110100100110: color_data = 12'b001111111111;
20'b00111101110100100111: color_data = 12'b001111111111;
20'b00111101110100101000: color_data = 12'b001111111111;
20'b00111101110100101001: color_data = 12'b001111111111;
20'b00111101110100101010: color_data = 12'b001111111111;
20'b00111101110100101011: color_data = 12'b001111111111;
20'b00111101110100101100: color_data = 12'b001111111111;
20'b00111101110100101101: color_data = 12'b001111111111;
20'b00111101110100101111: color_data = 12'b001111111111;
20'b00111101110100110000: color_data = 12'b001111111111;
20'b00111101110100110001: color_data = 12'b001111111111;
20'b00111101110100110010: color_data = 12'b001111111111;
20'b00111101110100110011: color_data = 12'b001111111111;
20'b00111101110100110100: color_data = 12'b001111111111;
20'b00111101110100110101: color_data = 12'b001111111111;
20'b00111101110100110110: color_data = 12'b001111111111;
20'b00111101110100110111: color_data = 12'b001111111111;
20'b00111101110100111000: color_data = 12'b001111111111;
20'b00111101110101000100: color_data = 12'b000011110111;
20'b00111101110101000101: color_data = 12'b000011110111;
20'b00111101110101000110: color_data = 12'b000011110111;
20'b00111101110101000111: color_data = 12'b000011110111;
20'b00111101110101001000: color_data = 12'b000011110111;
20'b00111101110101001001: color_data = 12'b000011110111;
20'b00111101110101001010: color_data = 12'b000011110111;
20'b00111101110101001011: color_data = 12'b000011110111;
20'b00111101110101001100: color_data = 12'b000011110111;
20'b00111101110101001101: color_data = 12'b000011110111;
20'b00111101110101001111: color_data = 12'b000011110111;
20'b00111101110101010000: color_data = 12'b000011110111;
20'b00111101110101010001: color_data = 12'b000011110111;
20'b00111101110101010010: color_data = 12'b000011110111;
20'b00111101110101010011: color_data = 12'b000011110111;
20'b00111101110101010100: color_data = 12'b000011110111;
20'b00111101110101010101: color_data = 12'b000011110111;
20'b00111101110101010110: color_data = 12'b000011110111;
20'b00111101110101010111: color_data = 12'b000011110111;
20'b00111101110101011000: color_data = 12'b000011110111;
20'b00111101110101011010: color_data = 12'b000011110111;
20'b00111101110101011011: color_data = 12'b000011110111;
20'b00111101110101011100: color_data = 12'b000011110111;
20'b00111101110101011101: color_data = 12'b000011110111;
20'b00111101110101011110: color_data = 12'b000011110111;
20'b00111101110101011111: color_data = 12'b000011110111;
20'b00111101110101100000: color_data = 12'b000011110111;
20'b00111101110101100001: color_data = 12'b000011110111;
20'b00111101110101100010: color_data = 12'b000011110111;
20'b00111101110101100011: color_data = 12'b000011110111;
20'b00111101110111010011: color_data = 12'b000000001111;
20'b00111101110111010100: color_data = 12'b000000001111;
20'b00111101110111010101: color_data = 12'b000000001111;
20'b00111101110111010110: color_data = 12'b000000001111;
20'b00111101110111010111: color_data = 12'b000000001111;
20'b00111101110111011000: color_data = 12'b000000001111;
20'b00111101110111011001: color_data = 12'b000000001111;
20'b00111101110111011010: color_data = 12'b000000001111;
20'b00111101110111011011: color_data = 12'b000000001111;
20'b00111101110111011100: color_data = 12'b000000001111;
20'b00111101110111011110: color_data = 12'b000000001111;
20'b00111101110111011111: color_data = 12'b000000001111;
20'b00111101110111100000: color_data = 12'b000000001111;
20'b00111101110111100001: color_data = 12'b000000001111;
20'b00111101110111100010: color_data = 12'b000000001111;
20'b00111101110111100011: color_data = 12'b000000001111;
20'b00111101110111100100: color_data = 12'b000000001111;
20'b00111101110111100101: color_data = 12'b000000001111;
20'b00111101110111100110: color_data = 12'b000000001111;
20'b00111101110111100111: color_data = 12'b000000001111;
20'b00111110000010100001: color_data = 12'b111100001111;
20'b00111110000010100010: color_data = 12'b111100001111;
20'b00111110000010100011: color_data = 12'b111100001111;
20'b00111110000010100100: color_data = 12'b111100001111;
20'b00111110000010100101: color_data = 12'b111100001111;
20'b00111110000010100110: color_data = 12'b111100001111;
20'b00111110000010100111: color_data = 12'b111100001111;
20'b00111110000010101000: color_data = 12'b111100001111;
20'b00111110000010101001: color_data = 12'b111100001111;
20'b00111110000010101010: color_data = 12'b111100001111;
20'b00111110000011101101: color_data = 12'b000001111111;
20'b00111110000011101110: color_data = 12'b000001111111;
20'b00111110000011101111: color_data = 12'b000001111111;
20'b00111110000011110000: color_data = 12'b000001111111;
20'b00111110000011110001: color_data = 12'b000001111111;
20'b00111110000011110010: color_data = 12'b000001111111;
20'b00111110000011110011: color_data = 12'b000001111111;
20'b00111110000011110100: color_data = 12'b000001111111;
20'b00111110000011110101: color_data = 12'b000001111111;
20'b00111110000011110110: color_data = 12'b000001111111;
20'b00111110000011111000: color_data = 12'b000001111111;
20'b00111110000011111001: color_data = 12'b000001111111;
20'b00111110000011111010: color_data = 12'b000001111111;
20'b00111110000011111011: color_data = 12'b000001111111;
20'b00111110000011111100: color_data = 12'b000001111111;
20'b00111110000011111101: color_data = 12'b000001111111;
20'b00111110000011111110: color_data = 12'b000001111111;
20'b00111110000011111111: color_data = 12'b000001111111;
20'b00111110000100000000: color_data = 12'b000001111111;
20'b00111110000100000001: color_data = 12'b000001111111;
20'b00111110000100100100: color_data = 12'b001111111111;
20'b00111110000100100101: color_data = 12'b001111111111;
20'b00111110000100100110: color_data = 12'b001111111111;
20'b00111110000100100111: color_data = 12'b001111111111;
20'b00111110000100101000: color_data = 12'b001111111111;
20'b00111110000100101001: color_data = 12'b001111111111;
20'b00111110000100101010: color_data = 12'b001111111111;
20'b00111110000100101011: color_data = 12'b001111111111;
20'b00111110000100101100: color_data = 12'b001111111111;
20'b00111110000100101101: color_data = 12'b001111111111;
20'b00111110000100101111: color_data = 12'b001111111111;
20'b00111110000100110000: color_data = 12'b001111111111;
20'b00111110000100110001: color_data = 12'b001111111111;
20'b00111110000100110010: color_data = 12'b001111111111;
20'b00111110000100110011: color_data = 12'b001111111111;
20'b00111110000100110100: color_data = 12'b001111111111;
20'b00111110000100110101: color_data = 12'b001111111111;
20'b00111110000100110110: color_data = 12'b001111111111;
20'b00111110000100110111: color_data = 12'b001111111111;
20'b00111110000100111000: color_data = 12'b001111111111;
20'b00111110000101000100: color_data = 12'b000011110111;
20'b00111110000101000101: color_data = 12'b000011110111;
20'b00111110000101000110: color_data = 12'b000011110111;
20'b00111110000101000111: color_data = 12'b000011110111;
20'b00111110000101001000: color_data = 12'b000011110111;
20'b00111110000101001001: color_data = 12'b000011110111;
20'b00111110000101001010: color_data = 12'b000011110111;
20'b00111110000101001011: color_data = 12'b000011110111;
20'b00111110000101001100: color_data = 12'b000011110111;
20'b00111110000101001101: color_data = 12'b000011110111;
20'b00111110000101001111: color_data = 12'b000011110111;
20'b00111110000101010000: color_data = 12'b000011110111;
20'b00111110000101010001: color_data = 12'b000011110111;
20'b00111110000101010010: color_data = 12'b000011110111;
20'b00111110000101010011: color_data = 12'b000011110111;
20'b00111110000101010100: color_data = 12'b000011110111;
20'b00111110000101010101: color_data = 12'b000011110111;
20'b00111110000101010110: color_data = 12'b000011110111;
20'b00111110000101010111: color_data = 12'b000011110111;
20'b00111110000101011000: color_data = 12'b000011110111;
20'b00111110000101011010: color_data = 12'b000011110111;
20'b00111110000101011011: color_data = 12'b000011110111;
20'b00111110000101011100: color_data = 12'b000011110111;
20'b00111110000101011101: color_data = 12'b000011110111;
20'b00111110000101011110: color_data = 12'b000011110111;
20'b00111110000101011111: color_data = 12'b000011110111;
20'b00111110000101100000: color_data = 12'b000011110111;
20'b00111110000101100001: color_data = 12'b000011110111;
20'b00111110000101100010: color_data = 12'b000011110111;
20'b00111110000101100011: color_data = 12'b000011110111;
20'b00111110000111010011: color_data = 12'b000000001111;
20'b00111110000111010100: color_data = 12'b000000001111;
20'b00111110000111010101: color_data = 12'b000000001111;
20'b00111110000111010110: color_data = 12'b000000001111;
20'b00111110000111010111: color_data = 12'b000000001111;
20'b00111110000111011000: color_data = 12'b000000001111;
20'b00111110000111011001: color_data = 12'b000000001111;
20'b00111110000111011010: color_data = 12'b000000001111;
20'b00111110000111011011: color_data = 12'b000000001111;
20'b00111110000111011100: color_data = 12'b000000001111;
20'b00111110000111011110: color_data = 12'b000000001111;
20'b00111110000111011111: color_data = 12'b000000001111;
20'b00111110000111100000: color_data = 12'b000000001111;
20'b00111110000111100001: color_data = 12'b000000001111;
20'b00111110000111100010: color_data = 12'b000000001111;
20'b00111110000111100011: color_data = 12'b000000001111;
20'b00111110000111100100: color_data = 12'b000000001111;
20'b00111110000111100101: color_data = 12'b000000001111;
20'b00111110000111100110: color_data = 12'b000000001111;
20'b00111110000111100111: color_data = 12'b000000001111;
20'b00111110010010100001: color_data = 12'b111100001111;
20'b00111110010010100010: color_data = 12'b111100001111;
20'b00111110010010100011: color_data = 12'b111100001111;
20'b00111110010010100100: color_data = 12'b111100001111;
20'b00111110010010100101: color_data = 12'b111100001111;
20'b00111110010010100110: color_data = 12'b111100001111;
20'b00111110010010100111: color_data = 12'b111100001111;
20'b00111110010010101000: color_data = 12'b111100001111;
20'b00111110010010101001: color_data = 12'b111100001111;
20'b00111110010010101010: color_data = 12'b111100001111;
20'b00111110010011101101: color_data = 12'b000001111111;
20'b00111110010011101110: color_data = 12'b000001111111;
20'b00111110010011101111: color_data = 12'b000001111111;
20'b00111110010011110000: color_data = 12'b000001111111;
20'b00111110010011110001: color_data = 12'b000001111111;
20'b00111110010011110010: color_data = 12'b000001111111;
20'b00111110010011110011: color_data = 12'b000001111111;
20'b00111110010011110100: color_data = 12'b000001111111;
20'b00111110010011110101: color_data = 12'b000001111111;
20'b00111110010011110110: color_data = 12'b000001111111;
20'b00111110010011111000: color_data = 12'b000001111111;
20'b00111110010011111001: color_data = 12'b000001111111;
20'b00111110010011111010: color_data = 12'b000001111111;
20'b00111110010011111011: color_data = 12'b000001111111;
20'b00111110010011111100: color_data = 12'b000001111111;
20'b00111110010011111101: color_data = 12'b000001111111;
20'b00111110010011111110: color_data = 12'b000001111111;
20'b00111110010011111111: color_data = 12'b000001111111;
20'b00111110010100000000: color_data = 12'b000001111111;
20'b00111110010100000001: color_data = 12'b000001111111;
20'b00111110010100100100: color_data = 12'b001111111111;
20'b00111110010100100101: color_data = 12'b001111111111;
20'b00111110010100100110: color_data = 12'b001111111111;
20'b00111110010100100111: color_data = 12'b001111111111;
20'b00111110010100101000: color_data = 12'b001111111111;
20'b00111110010100101001: color_data = 12'b001111111111;
20'b00111110010100101010: color_data = 12'b001111111111;
20'b00111110010100101011: color_data = 12'b001111111111;
20'b00111110010100101100: color_data = 12'b001111111111;
20'b00111110010100101101: color_data = 12'b001111111111;
20'b00111110010100101111: color_data = 12'b001111111111;
20'b00111110010100110000: color_data = 12'b001111111111;
20'b00111110010100110001: color_data = 12'b001111111111;
20'b00111110010100110010: color_data = 12'b001111111111;
20'b00111110010100110011: color_data = 12'b001111111111;
20'b00111110010100110100: color_data = 12'b001111111111;
20'b00111110010100110101: color_data = 12'b001111111111;
20'b00111110010100110110: color_data = 12'b001111111111;
20'b00111110010100110111: color_data = 12'b001111111111;
20'b00111110010100111000: color_data = 12'b001111111111;
20'b00111110010101000100: color_data = 12'b000011110111;
20'b00111110010101000101: color_data = 12'b000011110111;
20'b00111110010101000110: color_data = 12'b000011110111;
20'b00111110010101000111: color_data = 12'b000011110111;
20'b00111110010101001000: color_data = 12'b000011110111;
20'b00111110010101001001: color_data = 12'b000011110111;
20'b00111110010101001010: color_data = 12'b000011110111;
20'b00111110010101001011: color_data = 12'b000011110111;
20'b00111110010101001100: color_data = 12'b000011110111;
20'b00111110010101001101: color_data = 12'b000011110111;
20'b00111110010101001111: color_data = 12'b000011110111;
20'b00111110010101010000: color_data = 12'b000011110111;
20'b00111110010101010001: color_data = 12'b000011110111;
20'b00111110010101010010: color_data = 12'b000011110111;
20'b00111110010101010011: color_data = 12'b000011110111;
20'b00111110010101010100: color_data = 12'b000011110111;
20'b00111110010101010101: color_data = 12'b000011110111;
20'b00111110010101010110: color_data = 12'b000011110111;
20'b00111110010101010111: color_data = 12'b000011110111;
20'b00111110010101011000: color_data = 12'b000011110111;
20'b00111110010101011010: color_data = 12'b000011110111;
20'b00111110010101011011: color_data = 12'b000011110111;
20'b00111110010101011100: color_data = 12'b000011110111;
20'b00111110010101011101: color_data = 12'b000011110111;
20'b00111110010101011110: color_data = 12'b000011110111;
20'b00111110010101011111: color_data = 12'b000011110111;
20'b00111110010101100000: color_data = 12'b000011110111;
20'b00111110010101100001: color_data = 12'b000011110111;
20'b00111110010101100010: color_data = 12'b000011110111;
20'b00111110010101100011: color_data = 12'b000011110111;
20'b00111110010111010011: color_data = 12'b000000001111;
20'b00111110010111010100: color_data = 12'b000000001111;
20'b00111110010111010101: color_data = 12'b000000001111;
20'b00111110010111010110: color_data = 12'b000000001111;
20'b00111110010111010111: color_data = 12'b000000001111;
20'b00111110010111011000: color_data = 12'b000000001111;
20'b00111110010111011001: color_data = 12'b000000001111;
20'b00111110010111011010: color_data = 12'b000000001111;
20'b00111110010111011011: color_data = 12'b000000001111;
20'b00111110010111011100: color_data = 12'b000000001111;
20'b00111110010111011110: color_data = 12'b000000001111;
20'b00111110010111011111: color_data = 12'b000000001111;
20'b00111110010111100000: color_data = 12'b000000001111;
20'b00111110010111100001: color_data = 12'b000000001111;
20'b00111110010111100010: color_data = 12'b000000001111;
20'b00111110010111100011: color_data = 12'b000000001111;
20'b00111110010111100100: color_data = 12'b000000001111;
20'b00111110010111100101: color_data = 12'b000000001111;
20'b00111110010111100110: color_data = 12'b000000001111;
20'b00111110010111100111: color_data = 12'b000000001111;
20'b00111110100010100001: color_data = 12'b111100001111;
20'b00111110100010100010: color_data = 12'b111100001111;
20'b00111110100010100011: color_data = 12'b111100001111;
20'b00111110100010100100: color_data = 12'b111100001111;
20'b00111110100010100101: color_data = 12'b111100001111;
20'b00111110100010100110: color_data = 12'b111100001111;
20'b00111110100010100111: color_data = 12'b111100001111;
20'b00111110100010101000: color_data = 12'b111100001111;
20'b00111110100010101001: color_data = 12'b111100001111;
20'b00111110100010101010: color_data = 12'b111100001111;
20'b00111110100011101101: color_data = 12'b000001111111;
20'b00111110100011101110: color_data = 12'b000001111111;
20'b00111110100011101111: color_data = 12'b000001111111;
20'b00111110100011110000: color_data = 12'b000001111111;
20'b00111110100011110001: color_data = 12'b000001111111;
20'b00111110100011110010: color_data = 12'b000001111111;
20'b00111110100011110011: color_data = 12'b000001111111;
20'b00111110100011110100: color_data = 12'b000001111111;
20'b00111110100011110101: color_data = 12'b000001111111;
20'b00111110100011110110: color_data = 12'b000001111111;
20'b00111110100011111000: color_data = 12'b000001111111;
20'b00111110100011111001: color_data = 12'b000001111111;
20'b00111110100011111010: color_data = 12'b000001111111;
20'b00111110100011111011: color_data = 12'b000001111111;
20'b00111110100011111100: color_data = 12'b000001111111;
20'b00111110100011111101: color_data = 12'b000001111111;
20'b00111110100011111110: color_data = 12'b000001111111;
20'b00111110100011111111: color_data = 12'b000001111111;
20'b00111110100100000000: color_data = 12'b000001111111;
20'b00111110100100000001: color_data = 12'b000001111111;
20'b00111110100100100100: color_data = 12'b001111111111;
20'b00111110100100100101: color_data = 12'b001111111111;
20'b00111110100100100110: color_data = 12'b001111111111;
20'b00111110100100100111: color_data = 12'b001111111111;
20'b00111110100100101000: color_data = 12'b001111111111;
20'b00111110100100101001: color_data = 12'b001111111111;
20'b00111110100100101010: color_data = 12'b001111111111;
20'b00111110100100101011: color_data = 12'b001111111111;
20'b00111110100100101100: color_data = 12'b001111111111;
20'b00111110100100101101: color_data = 12'b001111111111;
20'b00111110100100101111: color_data = 12'b001111111111;
20'b00111110100100110000: color_data = 12'b001111111111;
20'b00111110100100110001: color_data = 12'b001111111111;
20'b00111110100100110010: color_data = 12'b001111111111;
20'b00111110100100110011: color_data = 12'b001111111111;
20'b00111110100100110100: color_data = 12'b001111111111;
20'b00111110100100110101: color_data = 12'b001111111111;
20'b00111110100100110110: color_data = 12'b001111111111;
20'b00111110100100110111: color_data = 12'b001111111111;
20'b00111110100100111000: color_data = 12'b001111111111;
20'b00111110100101000100: color_data = 12'b000011110111;
20'b00111110100101000101: color_data = 12'b000011110111;
20'b00111110100101000110: color_data = 12'b000011110111;
20'b00111110100101000111: color_data = 12'b000011110111;
20'b00111110100101001000: color_data = 12'b000011110111;
20'b00111110100101001001: color_data = 12'b000011110111;
20'b00111110100101001010: color_data = 12'b000011110111;
20'b00111110100101001011: color_data = 12'b000011110111;
20'b00111110100101001100: color_data = 12'b000011110111;
20'b00111110100101001101: color_data = 12'b000011110111;
20'b00111110100101001111: color_data = 12'b000011110111;
20'b00111110100101010000: color_data = 12'b000011110111;
20'b00111110100101010001: color_data = 12'b000011110111;
20'b00111110100101010010: color_data = 12'b000011110111;
20'b00111110100101010011: color_data = 12'b000011110111;
20'b00111110100101010100: color_data = 12'b000011110111;
20'b00111110100101010101: color_data = 12'b000011110111;
20'b00111110100101010110: color_data = 12'b000011110111;
20'b00111110100101010111: color_data = 12'b000011110111;
20'b00111110100101011000: color_data = 12'b000011110111;
20'b00111110100101011010: color_data = 12'b000011110111;
20'b00111110100101011011: color_data = 12'b000011110111;
20'b00111110100101011100: color_data = 12'b000011110111;
20'b00111110100101011101: color_data = 12'b000011110111;
20'b00111110100101011110: color_data = 12'b000011110111;
20'b00111110100101011111: color_data = 12'b000011110111;
20'b00111110100101100000: color_data = 12'b000011110111;
20'b00111110100101100001: color_data = 12'b000011110111;
20'b00111110100101100010: color_data = 12'b000011110111;
20'b00111110100101100011: color_data = 12'b000011110111;
20'b00111110100111010011: color_data = 12'b000000001111;
20'b00111110100111010100: color_data = 12'b000000001111;
20'b00111110100111010101: color_data = 12'b000000001111;
20'b00111110100111010110: color_data = 12'b000000001111;
20'b00111110100111010111: color_data = 12'b000000001111;
20'b00111110100111011000: color_data = 12'b000000001111;
20'b00111110100111011001: color_data = 12'b000000001111;
20'b00111110100111011010: color_data = 12'b000000001111;
20'b00111110100111011011: color_data = 12'b000000001111;
20'b00111110100111011100: color_data = 12'b000000001111;
20'b00111110100111011110: color_data = 12'b000000001111;
20'b00111110100111011111: color_data = 12'b000000001111;
20'b00111110100111100000: color_data = 12'b000000001111;
20'b00111110100111100001: color_data = 12'b000000001111;
20'b00111110100111100010: color_data = 12'b000000001111;
20'b00111110100111100011: color_data = 12'b000000001111;
20'b00111110100111100100: color_data = 12'b000000001111;
20'b00111110100111100101: color_data = 12'b000000001111;
20'b00111110100111100110: color_data = 12'b000000001111;
20'b00111110100111100111: color_data = 12'b000000001111;
20'b00111110110010100001: color_data = 12'b111100001111;
20'b00111110110010100010: color_data = 12'b111100001111;
20'b00111110110010100011: color_data = 12'b111100001111;
20'b00111110110010100100: color_data = 12'b111100001111;
20'b00111110110010100101: color_data = 12'b111100001111;
20'b00111110110010100110: color_data = 12'b111100001111;
20'b00111110110010100111: color_data = 12'b111100001111;
20'b00111110110010101000: color_data = 12'b111100001111;
20'b00111110110010101001: color_data = 12'b111100001111;
20'b00111110110010101010: color_data = 12'b111100001111;
20'b00111110110011101101: color_data = 12'b000001111111;
20'b00111110110011101110: color_data = 12'b000001111111;
20'b00111110110011101111: color_data = 12'b000001111111;
20'b00111110110011110000: color_data = 12'b000001111111;
20'b00111110110011110001: color_data = 12'b000001111111;
20'b00111110110011110010: color_data = 12'b000001111111;
20'b00111110110011110011: color_data = 12'b000001111111;
20'b00111110110011110100: color_data = 12'b000001111111;
20'b00111110110011110101: color_data = 12'b000001111111;
20'b00111110110011110110: color_data = 12'b000001111111;
20'b00111110110011111000: color_data = 12'b000001111111;
20'b00111110110011111001: color_data = 12'b000001111111;
20'b00111110110011111010: color_data = 12'b000001111111;
20'b00111110110011111011: color_data = 12'b000001111111;
20'b00111110110011111100: color_data = 12'b000001111111;
20'b00111110110011111101: color_data = 12'b000001111111;
20'b00111110110011111110: color_data = 12'b000001111111;
20'b00111110110011111111: color_data = 12'b000001111111;
20'b00111110110100000000: color_data = 12'b000001111111;
20'b00111110110100000001: color_data = 12'b000001111111;
20'b00111110110100100100: color_data = 12'b001111111111;
20'b00111110110100100101: color_data = 12'b001111111111;
20'b00111110110100100110: color_data = 12'b001111111111;
20'b00111110110100100111: color_data = 12'b001111111111;
20'b00111110110100101000: color_data = 12'b001111111111;
20'b00111110110100101001: color_data = 12'b001111111111;
20'b00111110110100101010: color_data = 12'b001111111111;
20'b00111110110100101011: color_data = 12'b001111111111;
20'b00111110110100101100: color_data = 12'b001111111111;
20'b00111110110100101101: color_data = 12'b001111111111;
20'b00111110110100101111: color_data = 12'b001111111111;
20'b00111110110100110000: color_data = 12'b001111111111;
20'b00111110110100110001: color_data = 12'b001111111111;
20'b00111110110100110010: color_data = 12'b001111111111;
20'b00111110110100110011: color_data = 12'b001111111111;
20'b00111110110100110100: color_data = 12'b001111111111;
20'b00111110110100110101: color_data = 12'b001111111111;
20'b00111110110100110110: color_data = 12'b001111111111;
20'b00111110110100110111: color_data = 12'b001111111111;
20'b00111110110100111000: color_data = 12'b001111111111;
20'b00111110110101000100: color_data = 12'b000011110111;
20'b00111110110101000101: color_data = 12'b000011110111;
20'b00111110110101000110: color_data = 12'b000011110111;
20'b00111110110101000111: color_data = 12'b000011110111;
20'b00111110110101001000: color_data = 12'b000011110111;
20'b00111110110101001001: color_data = 12'b000011110111;
20'b00111110110101001010: color_data = 12'b000011110111;
20'b00111110110101001011: color_data = 12'b000011110111;
20'b00111110110101001100: color_data = 12'b000011110111;
20'b00111110110101001101: color_data = 12'b000011110111;
20'b00111110110101001111: color_data = 12'b000011110111;
20'b00111110110101010000: color_data = 12'b000011110111;
20'b00111110110101010001: color_data = 12'b000011110111;
20'b00111110110101010010: color_data = 12'b000011110111;
20'b00111110110101010011: color_data = 12'b000011110111;
20'b00111110110101010100: color_data = 12'b000011110111;
20'b00111110110101010101: color_data = 12'b000011110111;
20'b00111110110101010110: color_data = 12'b000011110111;
20'b00111110110101010111: color_data = 12'b000011110111;
20'b00111110110101011000: color_data = 12'b000011110111;
20'b00111110110101011010: color_data = 12'b000011110111;
20'b00111110110101011011: color_data = 12'b000011110111;
20'b00111110110101011100: color_data = 12'b000011110111;
20'b00111110110101011101: color_data = 12'b000011110111;
20'b00111110110101011110: color_data = 12'b000011110111;
20'b00111110110101011111: color_data = 12'b000011110111;
20'b00111110110101100000: color_data = 12'b000011110111;
20'b00111110110101100001: color_data = 12'b000011110111;
20'b00111110110101100010: color_data = 12'b000011110111;
20'b00111110110101100011: color_data = 12'b000011110111;
20'b00111110110111010011: color_data = 12'b000000001111;
20'b00111110110111010100: color_data = 12'b000000001111;
20'b00111110110111010101: color_data = 12'b000000001111;
20'b00111110110111010110: color_data = 12'b000000001111;
20'b00111110110111010111: color_data = 12'b000000001111;
20'b00111110110111011000: color_data = 12'b000000001111;
20'b00111110110111011001: color_data = 12'b000000001111;
20'b00111110110111011010: color_data = 12'b000000001111;
20'b00111110110111011011: color_data = 12'b000000001111;
20'b00111110110111011100: color_data = 12'b000000001111;
20'b00111110110111011110: color_data = 12'b000000001111;
20'b00111110110111011111: color_data = 12'b000000001111;
20'b00111110110111100000: color_data = 12'b000000001111;
20'b00111110110111100001: color_data = 12'b000000001111;
20'b00111110110111100010: color_data = 12'b000000001111;
20'b00111110110111100011: color_data = 12'b000000001111;
20'b00111110110111100100: color_data = 12'b000000001111;
20'b00111110110111100101: color_data = 12'b000000001111;
20'b00111110110111100110: color_data = 12'b000000001111;
20'b00111110110111100111: color_data = 12'b000000001111;
20'b00111111000010100001: color_data = 12'b111100001111;
20'b00111111000010100010: color_data = 12'b111100001111;
20'b00111111000010100011: color_data = 12'b111100001111;
20'b00111111000010100100: color_data = 12'b111100001111;
20'b00111111000010100101: color_data = 12'b111100001111;
20'b00111111000010100110: color_data = 12'b111100001111;
20'b00111111000010100111: color_data = 12'b111100001111;
20'b00111111000010101000: color_data = 12'b111100001111;
20'b00111111000010101001: color_data = 12'b111100001111;
20'b00111111000010101010: color_data = 12'b111100001111;
20'b00111111000011101101: color_data = 12'b000001111111;
20'b00111111000011101110: color_data = 12'b000001111111;
20'b00111111000011101111: color_data = 12'b000001111111;
20'b00111111000011110000: color_data = 12'b000001111111;
20'b00111111000011110001: color_data = 12'b000001111111;
20'b00111111000011110010: color_data = 12'b000001111111;
20'b00111111000011110011: color_data = 12'b000001111111;
20'b00111111000011110100: color_data = 12'b000001111111;
20'b00111111000011110101: color_data = 12'b000001111111;
20'b00111111000011110110: color_data = 12'b000001111111;
20'b00111111000011111000: color_data = 12'b000001111111;
20'b00111111000011111001: color_data = 12'b000001111111;
20'b00111111000011111010: color_data = 12'b000001111111;
20'b00111111000011111011: color_data = 12'b000001111111;
20'b00111111000011111100: color_data = 12'b000001111111;
20'b00111111000011111101: color_data = 12'b000001111111;
20'b00111111000011111110: color_data = 12'b000001111111;
20'b00111111000011111111: color_data = 12'b000001111111;
20'b00111111000100000000: color_data = 12'b000001111111;
20'b00111111000100000001: color_data = 12'b000001111111;
20'b00111111000100100100: color_data = 12'b001111111111;
20'b00111111000100100101: color_data = 12'b001111111111;
20'b00111111000100100110: color_data = 12'b001111111111;
20'b00111111000100100111: color_data = 12'b001111111111;
20'b00111111000100101000: color_data = 12'b001111111111;
20'b00111111000100101001: color_data = 12'b001111111111;
20'b00111111000100101010: color_data = 12'b001111111111;
20'b00111111000100101011: color_data = 12'b001111111111;
20'b00111111000100101100: color_data = 12'b001111111111;
20'b00111111000100101101: color_data = 12'b001111111111;
20'b00111111000100101111: color_data = 12'b001111111111;
20'b00111111000100110000: color_data = 12'b001111111111;
20'b00111111000100110001: color_data = 12'b001111111111;
20'b00111111000100110010: color_data = 12'b001111111111;
20'b00111111000100110011: color_data = 12'b001111111111;
20'b00111111000100110100: color_data = 12'b001111111111;
20'b00111111000100110101: color_data = 12'b001111111111;
20'b00111111000100110110: color_data = 12'b001111111111;
20'b00111111000100110111: color_data = 12'b001111111111;
20'b00111111000100111000: color_data = 12'b001111111111;
20'b00111111000101000100: color_data = 12'b000011110111;
20'b00111111000101000101: color_data = 12'b000011110111;
20'b00111111000101000110: color_data = 12'b000011110111;
20'b00111111000101000111: color_data = 12'b000011110111;
20'b00111111000101001000: color_data = 12'b000011110111;
20'b00111111000101001001: color_data = 12'b000011110111;
20'b00111111000101001010: color_data = 12'b000011110111;
20'b00111111000101001011: color_data = 12'b000011110111;
20'b00111111000101001100: color_data = 12'b000011110111;
20'b00111111000101001101: color_data = 12'b000011110111;
20'b00111111000101001111: color_data = 12'b000011110111;
20'b00111111000101010000: color_data = 12'b000011110111;
20'b00111111000101010001: color_data = 12'b000011110111;
20'b00111111000101010010: color_data = 12'b000011110111;
20'b00111111000101010011: color_data = 12'b000011110111;
20'b00111111000101010100: color_data = 12'b000011110111;
20'b00111111000101010101: color_data = 12'b000011110111;
20'b00111111000101010110: color_data = 12'b000011110111;
20'b00111111000101010111: color_data = 12'b000011110111;
20'b00111111000101011000: color_data = 12'b000011110111;
20'b00111111000101011010: color_data = 12'b000011110111;
20'b00111111000101011011: color_data = 12'b000011110111;
20'b00111111000101011100: color_data = 12'b000011110111;
20'b00111111000101011101: color_data = 12'b000011110111;
20'b00111111000101011110: color_data = 12'b000011110111;
20'b00111111000101011111: color_data = 12'b000011110111;
20'b00111111000101100000: color_data = 12'b000011110111;
20'b00111111000101100001: color_data = 12'b000011110111;
20'b00111111000101100010: color_data = 12'b000011110111;
20'b00111111000101100011: color_data = 12'b000011110111;
20'b00111111000111010011: color_data = 12'b000000001111;
20'b00111111000111010100: color_data = 12'b000000001111;
20'b00111111000111010101: color_data = 12'b000000001111;
20'b00111111000111010110: color_data = 12'b000000001111;
20'b00111111000111010111: color_data = 12'b000000001111;
20'b00111111000111011000: color_data = 12'b000000001111;
20'b00111111000111011001: color_data = 12'b000000001111;
20'b00111111000111011010: color_data = 12'b000000001111;
20'b00111111000111011011: color_data = 12'b000000001111;
20'b00111111000111011100: color_data = 12'b000000001111;
20'b00111111000111011110: color_data = 12'b000000001111;
20'b00111111000111011111: color_data = 12'b000000001111;
20'b00111111000111100000: color_data = 12'b000000001111;
20'b00111111000111100001: color_data = 12'b000000001111;
20'b00111111000111100010: color_data = 12'b000000001111;
20'b00111111000111100011: color_data = 12'b000000001111;
20'b00111111000111100100: color_data = 12'b000000001111;
20'b00111111000111100101: color_data = 12'b000000001111;
20'b00111111000111100110: color_data = 12'b000000001111;
20'b00111111000111100111: color_data = 12'b000000001111;
20'b00111111010010100001: color_data = 12'b111100001111;
20'b00111111010010100010: color_data = 12'b111100001111;
20'b00111111010010100011: color_data = 12'b111100001111;
20'b00111111010010100100: color_data = 12'b111100001111;
20'b00111111010010100101: color_data = 12'b111100001111;
20'b00111111010010100110: color_data = 12'b111100001111;
20'b00111111010010100111: color_data = 12'b111100001111;
20'b00111111010010101000: color_data = 12'b111100001111;
20'b00111111010010101001: color_data = 12'b111100001111;
20'b00111111010010101010: color_data = 12'b111100001111;
20'b00111111010011101101: color_data = 12'b000001111111;
20'b00111111010011101110: color_data = 12'b000001111111;
20'b00111111010011101111: color_data = 12'b000001111111;
20'b00111111010011110000: color_data = 12'b000001111111;
20'b00111111010011110001: color_data = 12'b000001111111;
20'b00111111010011110010: color_data = 12'b000001111111;
20'b00111111010011110011: color_data = 12'b000001111111;
20'b00111111010011110100: color_data = 12'b000001111111;
20'b00111111010011110101: color_data = 12'b000001111111;
20'b00111111010011110110: color_data = 12'b000001111111;
20'b00111111010011111000: color_data = 12'b000001111111;
20'b00111111010011111001: color_data = 12'b000001111111;
20'b00111111010011111010: color_data = 12'b000001111111;
20'b00111111010011111011: color_data = 12'b000001111111;
20'b00111111010011111100: color_data = 12'b000001111111;
20'b00111111010011111101: color_data = 12'b000001111111;
20'b00111111010011111110: color_data = 12'b000001111111;
20'b00111111010011111111: color_data = 12'b000001111111;
20'b00111111010100000000: color_data = 12'b000001111111;
20'b00111111010100000001: color_data = 12'b000001111111;
20'b00111111010100100100: color_data = 12'b001111111111;
20'b00111111010100100101: color_data = 12'b001111111111;
20'b00111111010100100110: color_data = 12'b001111111111;
20'b00111111010100100111: color_data = 12'b001111111111;
20'b00111111010100101000: color_data = 12'b001111111111;
20'b00111111010100101001: color_data = 12'b001111111111;
20'b00111111010100101010: color_data = 12'b001111111111;
20'b00111111010100101011: color_data = 12'b001111111111;
20'b00111111010100101100: color_data = 12'b001111111111;
20'b00111111010100101101: color_data = 12'b001111111111;
20'b00111111010100101111: color_data = 12'b001111111111;
20'b00111111010100110000: color_data = 12'b001111111111;
20'b00111111010100110001: color_data = 12'b001111111111;
20'b00111111010100110010: color_data = 12'b001111111111;
20'b00111111010100110011: color_data = 12'b001111111111;
20'b00111111010100110100: color_data = 12'b001111111111;
20'b00111111010100110101: color_data = 12'b001111111111;
20'b00111111010100110110: color_data = 12'b001111111111;
20'b00111111010100110111: color_data = 12'b001111111111;
20'b00111111010100111000: color_data = 12'b001111111111;
20'b00111111010101000100: color_data = 12'b000011110111;
20'b00111111010101000101: color_data = 12'b000011110111;
20'b00111111010101000110: color_data = 12'b000011110111;
20'b00111111010101000111: color_data = 12'b000011110111;
20'b00111111010101001000: color_data = 12'b000011110111;
20'b00111111010101001001: color_data = 12'b000011110111;
20'b00111111010101001010: color_data = 12'b000011110111;
20'b00111111010101001011: color_data = 12'b000011110111;
20'b00111111010101001100: color_data = 12'b000011110111;
20'b00111111010101001101: color_data = 12'b000011110111;
20'b00111111010101001111: color_data = 12'b000011110111;
20'b00111111010101010000: color_data = 12'b000011110111;
20'b00111111010101010001: color_data = 12'b000011110111;
20'b00111111010101010010: color_data = 12'b000011110111;
20'b00111111010101010011: color_data = 12'b000011110111;
20'b00111111010101010100: color_data = 12'b000011110111;
20'b00111111010101010101: color_data = 12'b000011110111;
20'b00111111010101010110: color_data = 12'b000011110111;
20'b00111111010101010111: color_data = 12'b000011110111;
20'b00111111010101011000: color_data = 12'b000011110111;
20'b00111111010101011010: color_data = 12'b000011110111;
20'b00111111010101011011: color_data = 12'b000011110111;
20'b00111111010101011100: color_data = 12'b000011110111;
20'b00111111010101011101: color_data = 12'b000011110111;
20'b00111111010101011110: color_data = 12'b000011110111;
20'b00111111010101011111: color_data = 12'b000011110111;
20'b00111111010101100000: color_data = 12'b000011110111;
20'b00111111010101100001: color_data = 12'b000011110111;
20'b00111111010101100010: color_data = 12'b000011110111;
20'b00111111010101100011: color_data = 12'b000011110111;
20'b00111111010111010011: color_data = 12'b000000001111;
20'b00111111010111010100: color_data = 12'b000000001111;
20'b00111111010111010101: color_data = 12'b000000001111;
20'b00111111010111010110: color_data = 12'b000000001111;
20'b00111111010111010111: color_data = 12'b000000001111;
20'b00111111010111011000: color_data = 12'b000000001111;
20'b00111111010111011001: color_data = 12'b000000001111;
20'b00111111010111011010: color_data = 12'b000000001111;
20'b00111111010111011011: color_data = 12'b000000001111;
20'b00111111010111011100: color_data = 12'b000000001111;
20'b00111111010111011110: color_data = 12'b000000001111;
20'b00111111010111011111: color_data = 12'b000000001111;
20'b00111111010111100000: color_data = 12'b000000001111;
20'b00111111010111100001: color_data = 12'b000000001111;
20'b00111111010111100010: color_data = 12'b000000001111;
20'b00111111010111100011: color_data = 12'b000000001111;
20'b00111111010111100100: color_data = 12'b000000001111;
20'b00111111010111100101: color_data = 12'b000000001111;
20'b00111111010111100110: color_data = 12'b000000001111;
20'b00111111010111100111: color_data = 12'b000000001111;
20'b00111111100010100001: color_data = 12'b111100001111;
20'b00111111100010100010: color_data = 12'b111100001111;
20'b00111111100010100011: color_data = 12'b111100001111;
20'b00111111100010100100: color_data = 12'b111100001111;
20'b00111111100010100101: color_data = 12'b111100001111;
20'b00111111100010100110: color_data = 12'b111100001111;
20'b00111111100010100111: color_data = 12'b111100001111;
20'b00111111100010101000: color_data = 12'b111100001111;
20'b00111111100010101001: color_data = 12'b111100001111;
20'b00111111100010101010: color_data = 12'b111100001111;
20'b00111111100011101101: color_data = 12'b000001111111;
20'b00111111100011101110: color_data = 12'b000001111111;
20'b00111111100011101111: color_data = 12'b000001111111;
20'b00111111100011110000: color_data = 12'b000001111111;
20'b00111111100011110001: color_data = 12'b000001111111;
20'b00111111100011110010: color_data = 12'b000001111111;
20'b00111111100011110011: color_data = 12'b000001111111;
20'b00111111100011110100: color_data = 12'b000001111111;
20'b00111111100011110101: color_data = 12'b000001111111;
20'b00111111100011110110: color_data = 12'b000001111111;
20'b00111111100011111000: color_data = 12'b000001111111;
20'b00111111100011111001: color_data = 12'b000001111111;
20'b00111111100011111010: color_data = 12'b000001111111;
20'b00111111100011111011: color_data = 12'b000001111111;
20'b00111111100011111100: color_data = 12'b000001111111;
20'b00111111100011111101: color_data = 12'b000001111111;
20'b00111111100011111110: color_data = 12'b000001111111;
20'b00111111100011111111: color_data = 12'b000001111111;
20'b00111111100100000000: color_data = 12'b000001111111;
20'b00111111100100000001: color_data = 12'b000001111111;
20'b00111111100100100100: color_data = 12'b001111111111;
20'b00111111100100100101: color_data = 12'b001111111111;
20'b00111111100100100110: color_data = 12'b001111111111;
20'b00111111100100100111: color_data = 12'b001111111111;
20'b00111111100100101000: color_data = 12'b001111111111;
20'b00111111100100101001: color_data = 12'b001111111111;
20'b00111111100100101010: color_data = 12'b001111111111;
20'b00111111100100101011: color_data = 12'b001111111111;
20'b00111111100100101100: color_data = 12'b001111111111;
20'b00111111100100101101: color_data = 12'b001111111111;
20'b00111111100100101111: color_data = 12'b001111111111;
20'b00111111100100110000: color_data = 12'b001111111111;
20'b00111111100100110001: color_data = 12'b001111111111;
20'b00111111100100110010: color_data = 12'b001111111111;
20'b00111111100100110011: color_data = 12'b001111111111;
20'b00111111100100110100: color_data = 12'b001111111111;
20'b00111111100100110101: color_data = 12'b001111111111;
20'b00111111100100110110: color_data = 12'b001111111111;
20'b00111111100100110111: color_data = 12'b001111111111;
20'b00111111100100111000: color_data = 12'b001111111111;
20'b00111111100101000100: color_data = 12'b000011110111;
20'b00111111100101000101: color_data = 12'b000011110111;
20'b00111111100101000110: color_data = 12'b000011110111;
20'b00111111100101000111: color_data = 12'b000011110111;
20'b00111111100101001000: color_data = 12'b000011110111;
20'b00111111100101001001: color_data = 12'b000011110111;
20'b00111111100101001010: color_data = 12'b000011110111;
20'b00111111100101001011: color_data = 12'b000011110111;
20'b00111111100101001100: color_data = 12'b000011110111;
20'b00111111100101001101: color_data = 12'b000011110111;
20'b00111111100101001111: color_data = 12'b000011110111;
20'b00111111100101010000: color_data = 12'b000011110111;
20'b00111111100101010001: color_data = 12'b000011110111;
20'b00111111100101010010: color_data = 12'b000011110111;
20'b00111111100101010011: color_data = 12'b000011110111;
20'b00111111100101010100: color_data = 12'b000011110111;
20'b00111111100101010101: color_data = 12'b000011110111;
20'b00111111100101010110: color_data = 12'b000011110111;
20'b00111111100101010111: color_data = 12'b000011110111;
20'b00111111100101011000: color_data = 12'b000011110111;
20'b00111111100101011010: color_data = 12'b000011110111;
20'b00111111100101011011: color_data = 12'b000011110111;
20'b00111111100101011100: color_data = 12'b000011110111;
20'b00111111100101011101: color_data = 12'b000011110111;
20'b00111111100101011110: color_data = 12'b000011110111;
20'b00111111100101011111: color_data = 12'b000011110111;
20'b00111111100101100000: color_data = 12'b000011110111;
20'b00111111100101100001: color_data = 12'b000011110111;
20'b00111111100101100010: color_data = 12'b000011110111;
20'b00111111100101100011: color_data = 12'b000011110111;
20'b00111111100111010011: color_data = 12'b000000001111;
20'b00111111100111010100: color_data = 12'b000000001111;
20'b00111111100111010101: color_data = 12'b000000001111;
20'b00111111100111010110: color_data = 12'b000000001111;
20'b00111111100111010111: color_data = 12'b000000001111;
20'b00111111100111011000: color_data = 12'b000000001111;
20'b00111111100111011001: color_data = 12'b000000001111;
20'b00111111100111011010: color_data = 12'b000000001111;
20'b00111111100111011011: color_data = 12'b000000001111;
20'b00111111100111011100: color_data = 12'b000000001111;
20'b00111111100111011110: color_data = 12'b000000001111;
20'b00111111100111011111: color_data = 12'b000000001111;
20'b00111111100111100000: color_data = 12'b000000001111;
20'b00111111100111100001: color_data = 12'b000000001111;
20'b00111111100111100010: color_data = 12'b000000001111;
20'b00111111100111100011: color_data = 12'b000000001111;
20'b00111111100111100100: color_data = 12'b000000001111;
20'b00111111100111100101: color_data = 12'b000000001111;
20'b00111111100111100110: color_data = 12'b000000001111;
20'b00111111100111100111: color_data = 12'b000000001111;
20'b01000000000010110111: color_data = 12'b111011101110;
20'b01000000000010111000: color_data = 12'b111011101110;
20'b01000000000010111001: color_data = 12'b111011101110;
20'b01000000000010111010: color_data = 12'b111011101110;
20'b01000000000010111011: color_data = 12'b111011101110;
20'b01000000000010111100: color_data = 12'b111011101110;
20'b01000000000010111101: color_data = 12'b111011101110;
20'b01000000000010111110: color_data = 12'b111011101110;
20'b01000000000010111111: color_data = 12'b111011101110;
20'b01000000000011000000: color_data = 12'b111011101110;
20'b01000000000011000010: color_data = 12'b111011101110;
20'b01000000000011000011: color_data = 12'b111011101110;
20'b01000000000011000100: color_data = 12'b111011101110;
20'b01000000000011000101: color_data = 12'b111011101110;
20'b01000000000011000110: color_data = 12'b111011101110;
20'b01000000000011000111: color_data = 12'b111011101110;
20'b01000000000011001000: color_data = 12'b111011101110;
20'b01000000000011001001: color_data = 12'b111011101110;
20'b01000000000011001010: color_data = 12'b111011101110;
20'b01000000000011001011: color_data = 12'b111011101110;
20'b01000000000011001101: color_data = 12'b111011101110;
20'b01000000000011001110: color_data = 12'b111011101110;
20'b01000000000011001111: color_data = 12'b111011101110;
20'b01000000000011010000: color_data = 12'b111011101110;
20'b01000000000011010001: color_data = 12'b111011101110;
20'b01000000000011010010: color_data = 12'b111011101110;
20'b01000000000011010011: color_data = 12'b111011101110;
20'b01000000000011010100: color_data = 12'b111011101110;
20'b01000000000011010101: color_data = 12'b111011101110;
20'b01000000000011010110: color_data = 12'b111011101110;
20'b01000000000011111000: color_data = 12'b000001111111;
20'b01000000000011111001: color_data = 12'b000001111111;
20'b01000000000011111010: color_data = 12'b000001111111;
20'b01000000000011111011: color_data = 12'b000001111111;
20'b01000000000011111100: color_data = 12'b000001111111;
20'b01000000000011111101: color_data = 12'b000001111111;
20'b01000000000011111110: color_data = 12'b000001111111;
20'b01000000000011111111: color_data = 12'b000001111111;
20'b01000000000100000000: color_data = 12'b000001111111;
20'b01000000000100000001: color_data = 12'b000001111111;
20'b01000000000101000100: color_data = 12'b000011110111;
20'b01000000000101000101: color_data = 12'b000011110111;
20'b01000000000101000110: color_data = 12'b000011110111;
20'b01000000000101000111: color_data = 12'b000011110111;
20'b01000000000101001000: color_data = 12'b000011110111;
20'b01000000000101001001: color_data = 12'b000011110111;
20'b01000000000101001010: color_data = 12'b000011110111;
20'b01000000000101001011: color_data = 12'b000011110111;
20'b01000000000101001100: color_data = 12'b000011110111;
20'b01000000000101001101: color_data = 12'b000011110111;
20'b01000000000101100101: color_data = 12'b111011101110;
20'b01000000000101100110: color_data = 12'b111011101110;
20'b01000000000101100111: color_data = 12'b111011101110;
20'b01000000000101101000: color_data = 12'b111011101110;
20'b01000000000101101001: color_data = 12'b111011101110;
20'b01000000000101101010: color_data = 12'b111011101110;
20'b01000000000101101011: color_data = 12'b111011101110;
20'b01000000000101101100: color_data = 12'b111011101110;
20'b01000000000101101101: color_data = 12'b111011101110;
20'b01000000000101101110: color_data = 12'b111011101110;
20'b01000000000101110000: color_data = 12'b111011101110;
20'b01000000000101110001: color_data = 12'b111011101110;
20'b01000000000101110010: color_data = 12'b111011101110;
20'b01000000000101110011: color_data = 12'b111011101110;
20'b01000000000101110100: color_data = 12'b111011101110;
20'b01000000000101110101: color_data = 12'b111011101110;
20'b01000000000101110110: color_data = 12'b111011101110;
20'b01000000000101110111: color_data = 12'b111011101110;
20'b01000000000101111000: color_data = 12'b111011101110;
20'b01000000000101111001: color_data = 12'b111011101110;
20'b01000000000101111011: color_data = 12'b111011101110;
20'b01000000000101111100: color_data = 12'b111011101110;
20'b01000000000101111101: color_data = 12'b111011101110;
20'b01000000000101111110: color_data = 12'b111011101110;
20'b01000000000101111111: color_data = 12'b111011101110;
20'b01000000000110000000: color_data = 12'b111011101110;
20'b01000000000110000001: color_data = 12'b111011101110;
20'b01000000000110000010: color_data = 12'b111011101110;
20'b01000000000110000011: color_data = 12'b111011101110;
20'b01000000000110000100: color_data = 12'b111011101110;
20'b01000000000110000110: color_data = 12'b111011101110;
20'b01000000000110000111: color_data = 12'b111011101110;
20'b01000000000110001000: color_data = 12'b111011101110;
20'b01000000000110001001: color_data = 12'b111011101110;
20'b01000000000110001010: color_data = 12'b111011101110;
20'b01000000000110001011: color_data = 12'b111011101110;
20'b01000000000110001100: color_data = 12'b111011101110;
20'b01000000000110001101: color_data = 12'b111011101110;
20'b01000000000110001110: color_data = 12'b111011101110;
20'b01000000000110001111: color_data = 12'b111011101110;
20'b01000000000110100111: color_data = 12'b111011101110;
20'b01000000000110101000: color_data = 12'b111011101110;
20'b01000000000110101001: color_data = 12'b111011101110;
20'b01000000000110101010: color_data = 12'b111011101110;
20'b01000000000110101011: color_data = 12'b111011101110;
20'b01000000000110101100: color_data = 12'b111011101110;
20'b01000000000110101101: color_data = 12'b111011101110;
20'b01000000000110101110: color_data = 12'b111011101110;
20'b01000000000110101111: color_data = 12'b111011101110;
20'b01000000000110110000: color_data = 12'b111011101110;
20'b01000000000110110010: color_data = 12'b111011101110;
20'b01000000000110110011: color_data = 12'b111011101110;
20'b01000000000110110100: color_data = 12'b111011101110;
20'b01000000000110110101: color_data = 12'b111011101110;
20'b01000000000110110110: color_data = 12'b111011101110;
20'b01000000000110110111: color_data = 12'b111011101110;
20'b01000000000110111000: color_data = 12'b111011101110;
20'b01000000000110111001: color_data = 12'b111011101110;
20'b01000000000110111010: color_data = 12'b111011101110;
20'b01000000000110111011: color_data = 12'b111011101110;
20'b01000000000110111101: color_data = 12'b111011101110;
20'b01000000000110111110: color_data = 12'b111011101110;
20'b01000000000110111111: color_data = 12'b111011101110;
20'b01000000000111000000: color_data = 12'b111011101110;
20'b01000000000111000001: color_data = 12'b111011101110;
20'b01000000000111000010: color_data = 12'b111011101110;
20'b01000000000111000011: color_data = 12'b111011101110;
20'b01000000000111000100: color_data = 12'b111011101110;
20'b01000000000111000101: color_data = 12'b111011101110;
20'b01000000000111000110: color_data = 12'b111011101110;
20'b01000000000111001000: color_data = 12'b111011101110;
20'b01000000000111001001: color_data = 12'b111011101110;
20'b01000000000111001010: color_data = 12'b111011101110;
20'b01000000000111001011: color_data = 12'b111011101110;
20'b01000000000111001100: color_data = 12'b111011101110;
20'b01000000000111001101: color_data = 12'b111011101110;
20'b01000000000111001110: color_data = 12'b111011101110;
20'b01000000000111001111: color_data = 12'b111011101110;
20'b01000000000111010000: color_data = 12'b111011101110;
20'b01000000000111010001: color_data = 12'b111011101110;
20'b01000000010010110111: color_data = 12'b111011101110;
20'b01000000010010111000: color_data = 12'b111011101110;
20'b01000000010010111001: color_data = 12'b111011101110;
20'b01000000010010111010: color_data = 12'b111011101110;
20'b01000000010010111011: color_data = 12'b111011101110;
20'b01000000010010111100: color_data = 12'b111011101110;
20'b01000000010010111101: color_data = 12'b111011101110;
20'b01000000010010111110: color_data = 12'b111011101110;
20'b01000000010010111111: color_data = 12'b111011101110;
20'b01000000010011000000: color_data = 12'b111011101110;
20'b01000000010011000010: color_data = 12'b111011101110;
20'b01000000010011000011: color_data = 12'b111011101110;
20'b01000000010011000100: color_data = 12'b111011101110;
20'b01000000010011000101: color_data = 12'b111011101110;
20'b01000000010011000110: color_data = 12'b111011101110;
20'b01000000010011000111: color_data = 12'b111011101110;
20'b01000000010011001000: color_data = 12'b111011101110;
20'b01000000010011001001: color_data = 12'b111011101110;
20'b01000000010011001010: color_data = 12'b111011101110;
20'b01000000010011001011: color_data = 12'b111011101110;
20'b01000000010011001101: color_data = 12'b111011101110;
20'b01000000010011001110: color_data = 12'b111011101110;
20'b01000000010011001111: color_data = 12'b111011101110;
20'b01000000010011010000: color_data = 12'b111011101110;
20'b01000000010011010001: color_data = 12'b111011101110;
20'b01000000010011010010: color_data = 12'b111011101110;
20'b01000000010011010011: color_data = 12'b111011101110;
20'b01000000010011010100: color_data = 12'b111011101110;
20'b01000000010011010101: color_data = 12'b111011101110;
20'b01000000010011010110: color_data = 12'b111011101110;
20'b01000000010011111000: color_data = 12'b000001111111;
20'b01000000010011111001: color_data = 12'b000001111111;
20'b01000000010011111010: color_data = 12'b000001111111;
20'b01000000010011111011: color_data = 12'b000001111111;
20'b01000000010011111100: color_data = 12'b000001111111;
20'b01000000010011111101: color_data = 12'b000001111111;
20'b01000000010011111110: color_data = 12'b000001111111;
20'b01000000010011111111: color_data = 12'b000001111111;
20'b01000000010100000000: color_data = 12'b000001111111;
20'b01000000010100000001: color_data = 12'b000001111111;
20'b01000000010101000100: color_data = 12'b000011110111;
20'b01000000010101000101: color_data = 12'b000011110111;
20'b01000000010101000110: color_data = 12'b000011110111;
20'b01000000010101000111: color_data = 12'b000011110111;
20'b01000000010101001000: color_data = 12'b000011110111;
20'b01000000010101001001: color_data = 12'b000011110111;
20'b01000000010101001010: color_data = 12'b000011110111;
20'b01000000010101001011: color_data = 12'b000011110111;
20'b01000000010101001100: color_data = 12'b000011110111;
20'b01000000010101001101: color_data = 12'b000011110111;
20'b01000000010101100101: color_data = 12'b111011101110;
20'b01000000010101100110: color_data = 12'b111011101110;
20'b01000000010101100111: color_data = 12'b111011101110;
20'b01000000010101101000: color_data = 12'b111011101110;
20'b01000000010101101001: color_data = 12'b111011101110;
20'b01000000010101101010: color_data = 12'b111011101110;
20'b01000000010101101011: color_data = 12'b111011101110;
20'b01000000010101101100: color_data = 12'b111011101110;
20'b01000000010101101101: color_data = 12'b111011101110;
20'b01000000010101101110: color_data = 12'b111011101110;
20'b01000000010101110000: color_data = 12'b111011101110;
20'b01000000010101110001: color_data = 12'b111011101110;
20'b01000000010101110010: color_data = 12'b111011101110;
20'b01000000010101110011: color_data = 12'b111011101110;
20'b01000000010101110100: color_data = 12'b111011101110;
20'b01000000010101110101: color_data = 12'b111011101110;
20'b01000000010101110110: color_data = 12'b111011101110;
20'b01000000010101110111: color_data = 12'b111011101110;
20'b01000000010101111000: color_data = 12'b111011101110;
20'b01000000010101111001: color_data = 12'b111011101110;
20'b01000000010101111011: color_data = 12'b111011101110;
20'b01000000010101111100: color_data = 12'b111011101110;
20'b01000000010101111101: color_data = 12'b111011101110;
20'b01000000010101111110: color_data = 12'b111011101110;
20'b01000000010101111111: color_data = 12'b111011101110;
20'b01000000010110000000: color_data = 12'b111011101110;
20'b01000000010110000001: color_data = 12'b111011101110;
20'b01000000010110000010: color_data = 12'b111011101110;
20'b01000000010110000011: color_data = 12'b111011101110;
20'b01000000010110000100: color_data = 12'b111011101110;
20'b01000000010110000110: color_data = 12'b111011101110;
20'b01000000010110000111: color_data = 12'b111011101110;
20'b01000000010110001000: color_data = 12'b111011101110;
20'b01000000010110001001: color_data = 12'b111011101110;
20'b01000000010110001010: color_data = 12'b111011101110;
20'b01000000010110001011: color_data = 12'b111011101110;
20'b01000000010110001100: color_data = 12'b111011101110;
20'b01000000010110001101: color_data = 12'b111011101110;
20'b01000000010110001110: color_data = 12'b111011101110;
20'b01000000010110001111: color_data = 12'b111011101110;
20'b01000000010110100111: color_data = 12'b111011101110;
20'b01000000010110101000: color_data = 12'b111011101110;
20'b01000000010110101001: color_data = 12'b111011101110;
20'b01000000010110101010: color_data = 12'b111011101110;
20'b01000000010110101011: color_data = 12'b111011101110;
20'b01000000010110101100: color_data = 12'b111011101110;
20'b01000000010110101101: color_data = 12'b111011101110;
20'b01000000010110101110: color_data = 12'b111011101110;
20'b01000000010110101111: color_data = 12'b111011101110;
20'b01000000010110110000: color_data = 12'b111011101110;
20'b01000000010110110010: color_data = 12'b111011101110;
20'b01000000010110110011: color_data = 12'b111011101110;
20'b01000000010110110100: color_data = 12'b111011101110;
20'b01000000010110110101: color_data = 12'b111011101110;
20'b01000000010110110110: color_data = 12'b111011101110;
20'b01000000010110110111: color_data = 12'b111011101110;
20'b01000000010110111000: color_data = 12'b111011101110;
20'b01000000010110111001: color_data = 12'b111011101110;
20'b01000000010110111010: color_data = 12'b111011101110;
20'b01000000010110111011: color_data = 12'b111011101110;
20'b01000000010110111101: color_data = 12'b111011101110;
20'b01000000010110111110: color_data = 12'b111011101110;
20'b01000000010110111111: color_data = 12'b111011101110;
20'b01000000010111000000: color_data = 12'b111011101110;
20'b01000000010111000001: color_data = 12'b111011101110;
20'b01000000010111000010: color_data = 12'b111011101110;
20'b01000000010111000011: color_data = 12'b111011101110;
20'b01000000010111000100: color_data = 12'b111011101110;
20'b01000000010111000101: color_data = 12'b111011101110;
20'b01000000010111000110: color_data = 12'b111011101110;
20'b01000000010111001000: color_data = 12'b111011101110;
20'b01000000010111001001: color_data = 12'b111011101110;
20'b01000000010111001010: color_data = 12'b111011101110;
20'b01000000010111001011: color_data = 12'b111011101110;
20'b01000000010111001100: color_data = 12'b111011101110;
20'b01000000010111001101: color_data = 12'b111011101110;
20'b01000000010111001110: color_data = 12'b111011101110;
20'b01000000010111001111: color_data = 12'b111011101110;
20'b01000000010111010000: color_data = 12'b111011101110;
20'b01000000010111010001: color_data = 12'b111011101110;
20'b01000000100010110111: color_data = 12'b111011101110;
20'b01000000100010111000: color_data = 12'b111011101110;
20'b01000000100010111001: color_data = 12'b111011101110;
20'b01000000100010111010: color_data = 12'b111011101110;
20'b01000000100010111011: color_data = 12'b111011101110;
20'b01000000100010111100: color_data = 12'b111011101110;
20'b01000000100010111101: color_data = 12'b111011101110;
20'b01000000100010111110: color_data = 12'b111011101110;
20'b01000000100010111111: color_data = 12'b111011101110;
20'b01000000100011000000: color_data = 12'b111011101110;
20'b01000000100011000010: color_data = 12'b111011101110;
20'b01000000100011000011: color_data = 12'b111011101110;
20'b01000000100011000100: color_data = 12'b111011101110;
20'b01000000100011000101: color_data = 12'b111011101110;
20'b01000000100011000110: color_data = 12'b111011101110;
20'b01000000100011000111: color_data = 12'b111011101110;
20'b01000000100011001000: color_data = 12'b111011101110;
20'b01000000100011001001: color_data = 12'b111011101110;
20'b01000000100011001010: color_data = 12'b111011101110;
20'b01000000100011001011: color_data = 12'b111011101110;
20'b01000000100011001101: color_data = 12'b111011101110;
20'b01000000100011001110: color_data = 12'b111011101110;
20'b01000000100011001111: color_data = 12'b111011101110;
20'b01000000100011010000: color_data = 12'b111011101110;
20'b01000000100011010001: color_data = 12'b111011101110;
20'b01000000100011010010: color_data = 12'b111011101110;
20'b01000000100011010011: color_data = 12'b111011101110;
20'b01000000100011010100: color_data = 12'b111011101110;
20'b01000000100011010101: color_data = 12'b111011101110;
20'b01000000100011010110: color_data = 12'b111011101110;
20'b01000000100011111000: color_data = 12'b000001111111;
20'b01000000100011111001: color_data = 12'b000001111111;
20'b01000000100011111010: color_data = 12'b000001111111;
20'b01000000100011111011: color_data = 12'b000001111111;
20'b01000000100011111100: color_data = 12'b000001111111;
20'b01000000100011111101: color_data = 12'b000001111111;
20'b01000000100011111110: color_data = 12'b000001111111;
20'b01000000100011111111: color_data = 12'b000001111111;
20'b01000000100100000000: color_data = 12'b000001111111;
20'b01000000100100000001: color_data = 12'b000001111111;
20'b01000000100101000100: color_data = 12'b000011110111;
20'b01000000100101000101: color_data = 12'b000011110111;
20'b01000000100101000110: color_data = 12'b000011110111;
20'b01000000100101000111: color_data = 12'b000011110111;
20'b01000000100101001000: color_data = 12'b000011110111;
20'b01000000100101001001: color_data = 12'b000011110111;
20'b01000000100101001010: color_data = 12'b000011110111;
20'b01000000100101001011: color_data = 12'b000011110111;
20'b01000000100101001100: color_data = 12'b000011110111;
20'b01000000100101001101: color_data = 12'b000011110111;
20'b01000000100101100101: color_data = 12'b111011101110;
20'b01000000100101100110: color_data = 12'b111011101110;
20'b01000000100101100111: color_data = 12'b111011101110;
20'b01000000100101101000: color_data = 12'b111011101110;
20'b01000000100101101001: color_data = 12'b111011101110;
20'b01000000100101101010: color_data = 12'b111011101110;
20'b01000000100101101011: color_data = 12'b111011101110;
20'b01000000100101101100: color_data = 12'b111011101110;
20'b01000000100101101101: color_data = 12'b111011101110;
20'b01000000100101101110: color_data = 12'b111011101110;
20'b01000000100101110000: color_data = 12'b111011101110;
20'b01000000100101110001: color_data = 12'b111011101110;
20'b01000000100101110010: color_data = 12'b111011101110;
20'b01000000100101110011: color_data = 12'b111011101110;
20'b01000000100101110100: color_data = 12'b111011101110;
20'b01000000100101110101: color_data = 12'b111011101110;
20'b01000000100101110110: color_data = 12'b111011101110;
20'b01000000100101110111: color_data = 12'b111011101110;
20'b01000000100101111000: color_data = 12'b111011101110;
20'b01000000100101111001: color_data = 12'b111011101110;
20'b01000000100101111011: color_data = 12'b111011101110;
20'b01000000100101111100: color_data = 12'b111011101110;
20'b01000000100101111101: color_data = 12'b111011101110;
20'b01000000100101111110: color_data = 12'b111011101110;
20'b01000000100101111111: color_data = 12'b111011101110;
20'b01000000100110000000: color_data = 12'b111011101110;
20'b01000000100110000001: color_data = 12'b111011101110;
20'b01000000100110000010: color_data = 12'b111011101110;
20'b01000000100110000011: color_data = 12'b111011101110;
20'b01000000100110000100: color_data = 12'b111011101110;
20'b01000000100110000110: color_data = 12'b111011101110;
20'b01000000100110000111: color_data = 12'b111011101110;
20'b01000000100110001000: color_data = 12'b111011101110;
20'b01000000100110001001: color_data = 12'b111011101110;
20'b01000000100110001010: color_data = 12'b111011101110;
20'b01000000100110001011: color_data = 12'b111011101110;
20'b01000000100110001100: color_data = 12'b111011101110;
20'b01000000100110001101: color_data = 12'b111011101110;
20'b01000000100110001110: color_data = 12'b111011101110;
20'b01000000100110001111: color_data = 12'b111011101110;
20'b01000000100110100111: color_data = 12'b111011101110;
20'b01000000100110101000: color_data = 12'b111011101110;
20'b01000000100110101001: color_data = 12'b111011101110;
20'b01000000100110101010: color_data = 12'b111011101110;
20'b01000000100110101011: color_data = 12'b111011101110;
20'b01000000100110101100: color_data = 12'b111011101110;
20'b01000000100110101101: color_data = 12'b111011101110;
20'b01000000100110101110: color_data = 12'b111011101110;
20'b01000000100110101111: color_data = 12'b111011101110;
20'b01000000100110110000: color_data = 12'b111011101110;
20'b01000000100110110010: color_data = 12'b111011101110;
20'b01000000100110110011: color_data = 12'b111011101110;
20'b01000000100110110100: color_data = 12'b111011101110;
20'b01000000100110110101: color_data = 12'b111011101110;
20'b01000000100110110110: color_data = 12'b111011101110;
20'b01000000100110110111: color_data = 12'b111011101110;
20'b01000000100110111000: color_data = 12'b111011101110;
20'b01000000100110111001: color_data = 12'b111011101110;
20'b01000000100110111010: color_data = 12'b111011101110;
20'b01000000100110111011: color_data = 12'b111011101110;
20'b01000000100110111101: color_data = 12'b111011101110;
20'b01000000100110111110: color_data = 12'b111011101110;
20'b01000000100110111111: color_data = 12'b111011101110;
20'b01000000100111000000: color_data = 12'b111011101110;
20'b01000000100111000001: color_data = 12'b111011101110;
20'b01000000100111000010: color_data = 12'b111011101110;
20'b01000000100111000011: color_data = 12'b111011101110;
20'b01000000100111000100: color_data = 12'b111011101110;
20'b01000000100111000101: color_data = 12'b111011101110;
20'b01000000100111000110: color_data = 12'b111011101110;
20'b01000000100111001000: color_data = 12'b111011101110;
20'b01000000100111001001: color_data = 12'b111011101110;
20'b01000000100111001010: color_data = 12'b111011101110;
20'b01000000100111001011: color_data = 12'b111011101110;
20'b01000000100111001100: color_data = 12'b111011101110;
20'b01000000100111001101: color_data = 12'b111011101110;
20'b01000000100111001110: color_data = 12'b111011101110;
20'b01000000100111001111: color_data = 12'b111011101110;
20'b01000000100111010000: color_data = 12'b111011101110;
20'b01000000100111010001: color_data = 12'b111011101110;
20'b01000000110010110111: color_data = 12'b111011101110;
20'b01000000110010111000: color_data = 12'b111011101110;
20'b01000000110010111001: color_data = 12'b111011101110;
20'b01000000110010111010: color_data = 12'b111011101110;
20'b01000000110010111011: color_data = 12'b111011101110;
20'b01000000110010111100: color_data = 12'b111011101110;
20'b01000000110010111101: color_data = 12'b111011101110;
20'b01000000110010111110: color_data = 12'b111011101110;
20'b01000000110010111111: color_data = 12'b111011101110;
20'b01000000110011000000: color_data = 12'b111011101110;
20'b01000000110011000010: color_data = 12'b111011101110;
20'b01000000110011000011: color_data = 12'b111011101110;
20'b01000000110011000100: color_data = 12'b111011101110;
20'b01000000110011000101: color_data = 12'b111011101110;
20'b01000000110011000110: color_data = 12'b111011101110;
20'b01000000110011000111: color_data = 12'b111011101110;
20'b01000000110011001000: color_data = 12'b111011101110;
20'b01000000110011001001: color_data = 12'b111011101110;
20'b01000000110011001010: color_data = 12'b111011101110;
20'b01000000110011001011: color_data = 12'b111011101110;
20'b01000000110011001101: color_data = 12'b111011101110;
20'b01000000110011001110: color_data = 12'b111011101110;
20'b01000000110011001111: color_data = 12'b111011101110;
20'b01000000110011010000: color_data = 12'b111011101110;
20'b01000000110011010001: color_data = 12'b111011101110;
20'b01000000110011010010: color_data = 12'b111011101110;
20'b01000000110011010011: color_data = 12'b111011101110;
20'b01000000110011010100: color_data = 12'b111011101110;
20'b01000000110011010101: color_data = 12'b111011101110;
20'b01000000110011010110: color_data = 12'b111011101110;
20'b01000000110011111000: color_data = 12'b000001111111;
20'b01000000110011111001: color_data = 12'b000001111111;
20'b01000000110011111010: color_data = 12'b000001111111;
20'b01000000110011111011: color_data = 12'b000001111111;
20'b01000000110011111100: color_data = 12'b000001111111;
20'b01000000110011111101: color_data = 12'b000001111111;
20'b01000000110011111110: color_data = 12'b000001111111;
20'b01000000110011111111: color_data = 12'b000001111111;
20'b01000000110100000000: color_data = 12'b000001111111;
20'b01000000110100000001: color_data = 12'b000001111111;
20'b01000000110101000100: color_data = 12'b000011110111;
20'b01000000110101000101: color_data = 12'b000011110111;
20'b01000000110101000110: color_data = 12'b000011110111;
20'b01000000110101000111: color_data = 12'b000011110111;
20'b01000000110101001000: color_data = 12'b000011110111;
20'b01000000110101001001: color_data = 12'b000011110111;
20'b01000000110101001010: color_data = 12'b000011110111;
20'b01000000110101001011: color_data = 12'b000011110111;
20'b01000000110101001100: color_data = 12'b000011110111;
20'b01000000110101001101: color_data = 12'b000011110111;
20'b01000000110101100101: color_data = 12'b111011101110;
20'b01000000110101100110: color_data = 12'b111011101110;
20'b01000000110101100111: color_data = 12'b111011101110;
20'b01000000110101101000: color_data = 12'b111011101110;
20'b01000000110101101001: color_data = 12'b111011101110;
20'b01000000110101101010: color_data = 12'b111011101110;
20'b01000000110101101011: color_data = 12'b111011101110;
20'b01000000110101101100: color_data = 12'b111011101110;
20'b01000000110101101101: color_data = 12'b111011101110;
20'b01000000110101101110: color_data = 12'b111011101110;
20'b01000000110101110000: color_data = 12'b111011101110;
20'b01000000110101110001: color_data = 12'b111011101110;
20'b01000000110101110010: color_data = 12'b111011101110;
20'b01000000110101110011: color_data = 12'b111011101110;
20'b01000000110101110100: color_data = 12'b111011101110;
20'b01000000110101110101: color_data = 12'b111011101110;
20'b01000000110101110110: color_data = 12'b111011101110;
20'b01000000110101110111: color_data = 12'b111011101110;
20'b01000000110101111000: color_data = 12'b111011101110;
20'b01000000110101111001: color_data = 12'b111011101110;
20'b01000000110101111011: color_data = 12'b111011101110;
20'b01000000110101111100: color_data = 12'b111011101110;
20'b01000000110101111101: color_data = 12'b111011101110;
20'b01000000110101111110: color_data = 12'b111011101110;
20'b01000000110101111111: color_data = 12'b111011101110;
20'b01000000110110000000: color_data = 12'b111011101110;
20'b01000000110110000001: color_data = 12'b111011101110;
20'b01000000110110000010: color_data = 12'b111011101110;
20'b01000000110110000011: color_data = 12'b111011101110;
20'b01000000110110000100: color_data = 12'b111011101110;
20'b01000000110110000110: color_data = 12'b111011101110;
20'b01000000110110000111: color_data = 12'b111011101110;
20'b01000000110110001000: color_data = 12'b111011101110;
20'b01000000110110001001: color_data = 12'b111011101110;
20'b01000000110110001010: color_data = 12'b111011101110;
20'b01000000110110001011: color_data = 12'b111011101110;
20'b01000000110110001100: color_data = 12'b111011101110;
20'b01000000110110001101: color_data = 12'b111011101110;
20'b01000000110110001110: color_data = 12'b111011101110;
20'b01000000110110001111: color_data = 12'b111011101110;
20'b01000000110110100111: color_data = 12'b111011101110;
20'b01000000110110101000: color_data = 12'b111011101110;
20'b01000000110110101001: color_data = 12'b111011101110;
20'b01000000110110101010: color_data = 12'b111011101110;
20'b01000000110110101011: color_data = 12'b111011101110;
20'b01000000110110101100: color_data = 12'b111011101110;
20'b01000000110110101101: color_data = 12'b111011101110;
20'b01000000110110101110: color_data = 12'b111011101110;
20'b01000000110110101111: color_data = 12'b111011101110;
20'b01000000110110110000: color_data = 12'b111011101110;
20'b01000000110110110010: color_data = 12'b111011101110;
20'b01000000110110110011: color_data = 12'b111011101110;
20'b01000000110110110100: color_data = 12'b111011101110;
20'b01000000110110110101: color_data = 12'b111011101110;
20'b01000000110110110110: color_data = 12'b111011101110;
20'b01000000110110110111: color_data = 12'b111011101110;
20'b01000000110110111000: color_data = 12'b111011101110;
20'b01000000110110111001: color_data = 12'b111011101110;
20'b01000000110110111010: color_data = 12'b111011101110;
20'b01000000110110111011: color_data = 12'b111011101110;
20'b01000000110110111101: color_data = 12'b111011101110;
20'b01000000110110111110: color_data = 12'b111011101110;
20'b01000000110110111111: color_data = 12'b111011101110;
20'b01000000110111000000: color_data = 12'b111011101110;
20'b01000000110111000001: color_data = 12'b111011101110;
20'b01000000110111000010: color_data = 12'b111011101110;
20'b01000000110111000011: color_data = 12'b111011101110;
20'b01000000110111000100: color_data = 12'b111011101110;
20'b01000000110111000101: color_data = 12'b111011101110;
20'b01000000110111000110: color_data = 12'b111011101110;
20'b01000000110111001000: color_data = 12'b111011101110;
20'b01000000110111001001: color_data = 12'b111011101110;
20'b01000000110111001010: color_data = 12'b111011101110;
20'b01000000110111001011: color_data = 12'b111011101110;
20'b01000000110111001100: color_data = 12'b111011101110;
20'b01000000110111001101: color_data = 12'b111011101110;
20'b01000000110111001110: color_data = 12'b111011101110;
20'b01000000110111001111: color_data = 12'b111011101110;
20'b01000000110111010000: color_data = 12'b111011101110;
20'b01000000110111010001: color_data = 12'b111011101110;
20'b01000001000010110111: color_data = 12'b111011101110;
20'b01000001000010111000: color_data = 12'b111011101110;
20'b01000001000010111001: color_data = 12'b111011101110;
20'b01000001000010111010: color_data = 12'b111011101110;
20'b01000001000010111011: color_data = 12'b111011101110;
20'b01000001000010111100: color_data = 12'b111011101110;
20'b01000001000010111101: color_data = 12'b111011101110;
20'b01000001000010111110: color_data = 12'b111011101110;
20'b01000001000010111111: color_data = 12'b111011101110;
20'b01000001000011000000: color_data = 12'b111011101110;
20'b01000001000011000010: color_data = 12'b111011101110;
20'b01000001000011000011: color_data = 12'b111011101110;
20'b01000001000011000100: color_data = 12'b111011101110;
20'b01000001000011000101: color_data = 12'b111011101110;
20'b01000001000011000110: color_data = 12'b111011101110;
20'b01000001000011000111: color_data = 12'b111011101110;
20'b01000001000011001000: color_data = 12'b111011101110;
20'b01000001000011001001: color_data = 12'b111011101110;
20'b01000001000011001010: color_data = 12'b111011101110;
20'b01000001000011001011: color_data = 12'b111011101110;
20'b01000001000011001101: color_data = 12'b111011101110;
20'b01000001000011001110: color_data = 12'b111011101110;
20'b01000001000011001111: color_data = 12'b111011101110;
20'b01000001000011010000: color_data = 12'b111011101110;
20'b01000001000011010001: color_data = 12'b111011101110;
20'b01000001000011010010: color_data = 12'b111011101110;
20'b01000001000011010011: color_data = 12'b111011101110;
20'b01000001000011010100: color_data = 12'b111011101110;
20'b01000001000011010101: color_data = 12'b111011101110;
20'b01000001000011010110: color_data = 12'b111011101110;
20'b01000001000011111000: color_data = 12'b000001111111;
20'b01000001000011111001: color_data = 12'b000001111111;
20'b01000001000011111010: color_data = 12'b000001111111;
20'b01000001000011111011: color_data = 12'b000001111111;
20'b01000001000011111100: color_data = 12'b000001111111;
20'b01000001000011111101: color_data = 12'b000001111111;
20'b01000001000011111110: color_data = 12'b000001111111;
20'b01000001000011111111: color_data = 12'b000001111111;
20'b01000001000100000000: color_data = 12'b000001111111;
20'b01000001000100000001: color_data = 12'b000001111111;
20'b01000001000101000100: color_data = 12'b000011110111;
20'b01000001000101000101: color_data = 12'b000011110111;
20'b01000001000101000110: color_data = 12'b000011110111;
20'b01000001000101000111: color_data = 12'b000011110111;
20'b01000001000101001000: color_data = 12'b000011110111;
20'b01000001000101001001: color_data = 12'b000011110111;
20'b01000001000101001010: color_data = 12'b000011110111;
20'b01000001000101001011: color_data = 12'b000011110111;
20'b01000001000101001100: color_data = 12'b000011110111;
20'b01000001000101001101: color_data = 12'b000011110111;
20'b01000001000101100101: color_data = 12'b111011101110;
20'b01000001000101100110: color_data = 12'b111011101110;
20'b01000001000101100111: color_data = 12'b111011101110;
20'b01000001000101101000: color_data = 12'b111011101110;
20'b01000001000101101001: color_data = 12'b111011101110;
20'b01000001000101101010: color_data = 12'b111011101110;
20'b01000001000101101011: color_data = 12'b111011101110;
20'b01000001000101101100: color_data = 12'b111011101110;
20'b01000001000101101101: color_data = 12'b111011101110;
20'b01000001000101101110: color_data = 12'b111011101110;
20'b01000001000101110000: color_data = 12'b111011101110;
20'b01000001000101110001: color_data = 12'b111011101110;
20'b01000001000101110010: color_data = 12'b111011101110;
20'b01000001000101110011: color_data = 12'b111011101110;
20'b01000001000101110100: color_data = 12'b111011101110;
20'b01000001000101110101: color_data = 12'b111011101110;
20'b01000001000101110110: color_data = 12'b111011101110;
20'b01000001000101110111: color_data = 12'b111011101110;
20'b01000001000101111000: color_data = 12'b111011101110;
20'b01000001000101111001: color_data = 12'b111011101110;
20'b01000001000101111011: color_data = 12'b111011101110;
20'b01000001000101111100: color_data = 12'b111011101110;
20'b01000001000101111101: color_data = 12'b111011101110;
20'b01000001000101111110: color_data = 12'b111011101110;
20'b01000001000101111111: color_data = 12'b111011101110;
20'b01000001000110000000: color_data = 12'b111011101110;
20'b01000001000110000001: color_data = 12'b111011101110;
20'b01000001000110000010: color_data = 12'b111011101110;
20'b01000001000110000011: color_data = 12'b111011101110;
20'b01000001000110000100: color_data = 12'b111011101110;
20'b01000001000110000110: color_data = 12'b111011101110;
20'b01000001000110000111: color_data = 12'b111011101110;
20'b01000001000110001000: color_data = 12'b111011101110;
20'b01000001000110001001: color_data = 12'b111011101110;
20'b01000001000110001010: color_data = 12'b111011101110;
20'b01000001000110001011: color_data = 12'b111011101110;
20'b01000001000110001100: color_data = 12'b111011101110;
20'b01000001000110001101: color_data = 12'b111011101110;
20'b01000001000110001110: color_data = 12'b111011101110;
20'b01000001000110001111: color_data = 12'b111011101110;
20'b01000001000110100111: color_data = 12'b111011101110;
20'b01000001000110101000: color_data = 12'b111011101110;
20'b01000001000110101001: color_data = 12'b111011101110;
20'b01000001000110101010: color_data = 12'b111011101110;
20'b01000001000110101011: color_data = 12'b111011101110;
20'b01000001000110101100: color_data = 12'b111011101110;
20'b01000001000110101101: color_data = 12'b111011101110;
20'b01000001000110101110: color_data = 12'b111011101110;
20'b01000001000110101111: color_data = 12'b111011101110;
20'b01000001000110110000: color_data = 12'b111011101110;
20'b01000001000110110010: color_data = 12'b111011101110;
20'b01000001000110110011: color_data = 12'b111011101110;
20'b01000001000110110100: color_data = 12'b111011101110;
20'b01000001000110110101: color_data = 12'b111011101110;
20'b01000001000110110110: color_data = 12'b111011101110;
20'b01000001000110110111: color_data = 12'b111011101110;
20'b01000001000110111000: color_data = 12'b111011101110;
20'b01000001000110111001: color_data = 12'b111011101110;
20'b01000001000110111010: color_data = 12'b111011101110;
20'b01000001000110111011: color_data = 12'b111011101110;
20'b01000001000110111101: color_data = 12'b111011101110;
20'b01000001000110111110: color_data = 12'b111011101110;
20'b01000001000110111111: color_data = 12'b111011101110;
20'b01000001000111000000: color_data = 12'b111011101110;
20'b01000001000111000001: color_data = 12'b111011101110;
20'b01000001000111000010: color_data = 12'b111011101110;
20'b01000001000111000011: color_data = 12'b111011101110;
20'b01000001000111000100: color_data = 12'b111011101110;
20'b01000001000111000101: color_data = 12'b111011101110;
20'b01000001000111000110: color_data = 12'b111011101110;
20'b01000001000111001000: color_data = 12'b111011101110;
20'b01000001000111001001: color_data = 12'b111011101110;
20'b01000001000111001010: color_data = 12'b111011101110;
20'b01000001000111001011: color_data = 12'b111011101110;
20'b01000001000111001100: color_data = 12'b111011101110;
20'b01000001000111001101: color_data = 12'b111011101110;
20'b01000001000111001110: color_data = 12'b111011101110;
20'b01000001000111001111: color_data = 12'b111011101110;
20'b01000001000111010000: color_data = 12'b111011101110;
20'b01000001000111010001: color_data = 12'b111011101110;
20'b01000001010010110111: color_data = 12'b111011101110;
20'b01000001010010111000: color_data = 12'b111011101110;
20'b01000001010010111001: color_data = 12'b111011101110;
20'b01000001010010111010: color_data = 12'b111011101110;
20'b01000001010010111011: color_data = 12'b111011101110;
20'b01000001010010111100: color_data = 12'b111011101110;
20'b01000001010010111101: color_data = 12'b111011101110;
20'b01000001010010111110: color_data = 12'b111011101110;
20'b01000001010010111111: color_data = 12'b111011101110;
20'b01000001010011000000: color_data = 12'b111011101110;
20'b01000001010011000010: color_data = 12'b111011101110;
20'b01000001010011000011: color_data = 12'b111011101110;
20'b01000001010011000100: color_data = 12'b111011101110;
20'b01000001010011000101: color_data = 12'b111011101110;
20'b01000001010011000110: color_data = 12'b111011101110;
20'b01000001010011000111: color_data = 12'b111011101110;
20'b01000001010011001000: color_data = 12'b111011101110;
20'b01000001010011001001: color_data = 12'b111011101110;
20'b01000001010011001010: color_data = 12'b111011101110;
20'b01000001010011001011: color_data = 12'b111011101110;
20'b01000001010011001101: color_data = 12'b111011101110;
20'b01000001010011001110: color_data = 12'b111011101110;
20'b01000001010011001111: color_data = 12'b111011101110;
20'b01000001010011010000: color_data = 12'b111011101110;
20'b01000001010011010001: color_data = 12'b111011101110;
20'b01000001010011010010: color_data = 12'b111011101110;
20'b01000001010011010011: color_data = 12'b111011101110;
20'b01000001010011010100: color_data = 12'b111011101110;
20'b01000001010011010101: color_data = 12'b111011101110;
20'b01000001010011010110: color_data = 12'b111011101110;
20'b01000001010011111000: color_data = 12'b000001111111;
20'b01000001010011111001: color_data = 12'b000001111111;
20'b01000001010011111010: color_data = 12'b000001111111;
20'b01000001010011111011: color_data = 12'b000001111111;
20'b01000001010011111100: color_data = 12'b000001111111;
20'b01000001010011111101: color_data = 12'b000001111111;
20'b01000001010011111110: color_data = 12'b000001111111;
20'b01000001010011111111: color_data = 12'b000001111111;
20'b01000001010100000000: color_data = 12'b000001111111;
20'b01000001010100000001: color_data = 12'b000001111111;
20'b01000001010101000100: color_data = 12'b000011110111;
20'b01000001010101000101: color_data = 12'b000011110111;
20'b01000001010101000110: color_data = 12'b000011110111;
20'b01000001010101000111: color_data = 12'b000011110111;
20'b01000001010101001000: color_data = 12'b000011110111;
20'b01000001010101001001: color_data = 12'b000011110111;
20'b01000001010101001010: color_data = 12'b000011110111;
20'b01000001010101001011: color_data = 12'b000011110111;
20'b01000001010101001100: color_data = 12'b000011110111;
20'b01000001010101001101: color_data = 12'b000011110111;
20'b01000001010101100101: color_data = 12'b111011101110;
20'b01000001010101100110: color_data = 12'b111011101110;
20'b01000001010101100111: color_data = 12'b111011101110;
20'b01000001010101101000: color_data = 12'b111011101110;
20'b01000001010101101001: color_data = 12'b111011101110;
20'b01000001010101101010: color_data = 12'b111011101110;
20'b01000001010101101011: color_data = 12'b111011101110;
20'b01000001010101101100: color_data = 12'b111011101110;
20'b01000001010101101101: color_data = 12'b111011101110;
20'b01000001010101101110: color_data = 12'b111011101110;
20'b01000001010101110000: color_data = 12'b111011101110;
20'b01000001010101110001: color_data = 12'b111011101110;
20'b01000001010101110010: color_data = 12'b111011101110;
20'b01000001010101110011: color_data = 12'b111011101110;
20'b01000001010101110100: color_data = 12'b111011101110;
20'b01000001010101110101: color_data = 12'b111011101110;
20'b01000001010101110110: color_data = 12'b111011101110;
20'b01000001010101110111: color_data = 12'b111011101110;
20'b01000001010101111000: color_data = 12'b111011101110;
20'b01000001010101111001: color_data = 12'b111011101110;
20'b01000001010101111011: color_data = 12'b111011101110;
20'b01000001010101111100: color_data = 12'b111011101110;
20'b01000001010101111101: color_data = 12'b111011101110;
20'b01000001010101111110: color_data = 12'b111011101110;
20'b01000001010101111111: color_data = 12'b111011101110;
20'b01000001010110000000: color_data = 12'b111011101110;
20'b01000001010110000001: color_data = 12'b111011101110;
20'b01000001010110000010: color_data = 12'b111011101110;
20'b01000001010110000011: color_data = 12'b111011101110;
20'b01000001010110000100: color_data = 12'b111011101110;
20'b01000001010110000110: color_data = 12'b111011101110;
20'b01000001010110000111: color_data = 12'b111011101110;
20'b01000001010110001000: color_data = 12'b111011101110;
20'b01000001010110001001: color_data = 12'b111011101110;
20'b01000001010110001010: color_data = 12'b111011101110;
20'b01000001010110001011: color_data = 12'b111011101110;
20'b01000001010110001100: color_data = 12'b111011101110;
20'b01000001010110001101: color_data = 12'b111011101110;
20'b01000001010110001110: color_data = 12'b111011101110;
20'b01000001010110001111: color_data = 12'b111011101110;
20'b01000001010110100111: color_data = 12'b111011101110;
20'b01000001010110101000: color_data = 12'b111011101110;
20'b01000001010110101001: color_data = 12'b111011101110;
20'b01000001010110101010: color_data = 12'b111011101110;
20'b01000001010110101011: color_data = 12'b111011101110;
20'b01000001010110101100: color_data = 12'b111011101110;
20'b01000001010110101101: color_data = 12'b111011101110;
20'b01000001010110101110: color_data = 12'b111011101110;
20'b01000001010110101111: color_data = 12'b111011101110;
20'b01000001010110110000: color_data = 12'b111011101110;
20'b01000001010110110010: color_data = 12'b111011101110;
20'b01000001010110110011: color_data = 12'b111011101110;
20'b01000001010110110100: color_data = 12'b111011101110;
20'b01000001010110110101: color_data = 12'b111011101110;
20'b01000001010110110110: color_data = 12'b111011101110;
20'b01000001010110110111: color_data = 12'b111011101110;
20'b01000001010110111000: color_data = 12'b111011101110;
20'b01000001010110111001: color_data = 12'b111011101110;
20'b01000001010110111010: color_data = 12'b111011101110;
20'b01000001010110111011: color_data = 12'b111011101110;
20'b01000001010110111101: color_data = 12'b111011101110;
20'b01000001010110111110: color_data = 12'b111011101110;
20'b01000001010110111111: color_data = 12'b111011101110;
20'b01000001010111000000: color_data = 12'b111011101110;
20'b01000001010111000001: color_data = 12'b111011101110;
20'b01000001010111000010: color_data = 12'b111011101110;
20'b01000001010111000011: color_data = 12'b111011101110;
20'b01000001010111000100: color_data = 12'b111011101110;
20'b01000001010111000101: color_data = 12'b111011101110;
20'b01000001010111000110: color_data = 12'b111011101110;
20'b01000001010111001000: color_data = 12'b111011101110;
20'b01000001010111001001: color_data = 12'b111011101110;
20'b01000001010111001010: color_data = 12'b111011101110;
20'b01000001010111001011: color_data = 12'b111011101110;
20'b01000001010111001100: color_data = 12'b111011101110;
20'b01000001010111001101: color_data = 12'b111011101110;
20'b01000001010111001110: color_data = 12'b111011101110;
20'b01000001010111001111: color_data = 12'b111011101110;
20'b01000001010111010000: color_data = 12'b111011101110;
20'b01000001010111010001: color_data = 12'b111011101110;
20'b01000001100010110111: color_data = 12'b111011101110;
20'b01000001100010111000: color_data = 12'b111011101110;
20'b01000001100010111001: color_data = 12'b111011101110;
20'b01000001100010111010: color_data = 12'b111011101110;
20'b01000001100010111011: color_data = 12'b111011101110;
20'b01000001100010111100: color_data = 12'b111011101110;
20'b01000001100010111101: color_data = 12'b111011101110;
20'b01000001100010111110: color_data = 12'b111011101110;
20'b01000001100010111111: color_data = 12'b111011101110;
20'b01000001100011000000: color_data = 12'b111011101110;
20'b01000001100011000010: color_data = 12'b111011101110;
20'b01000001100011000011: color_data = 12'b111011101110;
20'b01000001100011000100: color_data = 12'b111011101110;
20'b01000001100011000101: color_data = 12'b111011101110;
20'b01000001100011000110: color_data = 12'b111011101110;
20'b01000001100011000111: color_data = 12'b111011101110;
20'b01000001100011001000: color_data = 12'b111011101110;
20'b01000001100011001001: color_data = 12'b111011101110;
20'b01000001100011001010: color_data = 12'b111011101110;
20'b01000001100011001011: color_data = 12'b111011101110;
20'b01000001100011001101: color_data = 12'b111011101110;
20'b01000001100011001110: color_data = 12'b111011101110;
20'b01000001100011001111: color_data = 12'b111011101110;
20'b01000001100011010000: color_data = 12'b111011101110;
20'b01000001100011010001: color_data = 12'b111011101110;
20'b01000001100011010010: color_data = 12'b111011101110;
20'b01000001100011010011: color_data = 12'b111011101110;
20'b01000001100011010100: color_data = 12'b111011101110;
20'b01000001100011010101: color_data = 12'b111011101110;
20'b01000001100011010110: color_data = 12'b111011101110;
20'b01000001100011111000: color_data = 12'b000001111111;
20'b01000001100011111001: color_data = 12'b000001111111;
20'b01000001100011111010: color_data = 12'b000001111111;
20'b01000001100011111011: color_data = 12'b000001111111;
20'b01000001100011111100: color_data = 12'b000001111111;
20'b01000001100011111101: color_data = 12'b000001111111;
20'b01000001100011111110: color_data = 12'b000001111111;
20'b01000001100011111111: color_data = 12'b000001111111;
20'b01000001100100000000: color_data = 12'b000001111111;
20'b01000001100100000001: color_data = 12'b000001111111;
20'b01000001100101000100: color_data = 12'b000011110111;
20'b01000001100101000101: color_data = 12'b000011110111;
20'b01000001100101000110: color_data = 12'b000011110111;
20'b01000001100101000111: color_data = 12'b000011110111;
20'b01000001100101001000: color_data = 12'b000011110111;
20'b01000001100101001001: color_data = 12'b000011110111;
20'b01000001100101001010: color_data = 12'b000011110111;
20'b01000001100101001011: color_data = 12'b000011110111;
20'b01000001100101001100: color_data = 12'b000011110111;
20'b01000001100101001101: color_data = 12'b000011110111;
20'b01000001100101100101: color_data = 12'b111011101110;
20'b01000001100101100110: color_data = 12'b111011101110;
20'b01000001100101100111: color_data = 12'b111011101110;
20'b01000001100101101000: color_data = 12'b111011101110;
20'b01000001100101101001: color_data = 12'b111011101110;
20'b01000001100101101010: color_data = 12'b111011101110;
20'b01000001100101101011: color_data = 12'b111011101110;
20'b01000001100101101100: color_data = 12'b111011101110;
20'b01000001100101101101: color_data = 12'b111011101110;
20'b01000001100101101110: color_data = 12'b111011101110;
20'b01000001100101110000: color_data = 12'b111011101110;
20'b01000001100101110001: color_data = 12'b111011101110;
20'b01000001100101110010: color_data = 12'b111011101110;
20'b01000001100101110011: color_data = 12'b111011101110;
20'b01000001100101110100: color_data = 12'b111011101110;
20'b01000001100101110101: color_data = 12'b111011101110;
20'b01000001100101110110: color_data = 12'b111011101110;
20'b01000001100101110111: color_data = 12'b111011101110;
20'b01000001100101111000: color_data = 12'b111011101110;
20'b01000001100101111001: color_data = 12'b111011101110;
20'b01000001100101111011: color_data = 12'b111011101110;
20'b01000001100101111100: color_data = 12'b111011101110;
20'b01000001100101111101: color_data = 12'b111011101110;
20'b01000001100101111110: color_data = 12'b111011101110;
20'b01000001100101111111: color_data = 12'b111011101110;
20'b01000001100110000000: color_data = 12'b111011101110;
20'b01000001100110000001: color_data = 12'b111011101110;
20'b01000001100110000010: color_data = 12'b111011101110;
20'b01000001100110000011: color_data = 12'b111011101110;
20'b01000001100110000100: color_data = 12'b111011101110;
20'b01000001100110000110: color_data = 12'b111011101110;
20'b01000001100110000111: color_data = 12'b111011101110;
20'b01000001100110001000: color_data = 12'b111011101110;
20'b01000001100110001001: color_data = 12'b111011101110;
20'b01000001100110001010: color_data = 12'b111011101110;
20'b01000001100110001011: color_data = 12'b111011101110;
20'b01000001100110001100: color_data = 12'b111011101110;
20'b01000001100110001101: color_data = 12'b111011101110;
20'b01000001100110001110: color_data = 12'b111011101110;
20'b01000001100110001111: color_data = 12'b111011101110;
20'b01000001100110100111: color_data = 12'b111011101110;
20'b01000001100110101000: color_data = 12'b111011101110;
20'b01000001100110101001: color_data = 12'b111011101110;
20'b01000001100110101010: color_data = 12'b111011101110;
20'b01000001100110101011: color_data = 12'b111011101110;
20'b01000001100110101100: color_data = 12'b111011101110;
20'b01000001100110101101: color_data = 12'b111011101110;
20'b01000001100110101110: color_data = 12'b111011101110;
20'b01000001100110101111: color_data = 12'b111011101110;
20'b01000001100110110000: color_data = 12'b111011101110;
20'b01000001100110110010: color_data = 12'b111011101110;
20'b01000001100110110011: color_data = 12'b111011101110;
20'b01000001100110110100: color_data = 12'b111011101110;
20'b01000001100110110101: color_data = 12'b111011101110;
20'b01000001100110110110: color_data = 12'b111011101110;
20'b01000001100110110111: color_data = 12'b111011101110;
20'b01000001100110111000: color_data = 12'b111011101110;
20'b01000001100110111001: color_data = 12'b111011101110;
20'b01000001100110111010: color_data = 12'b111011101110;
20'b01000001100110111011: color_data = 12'b111011101110;
20'b01000001100110111101: color_data = 12'b111011101110;
20'b01000001100110111110: color_data = 12'b111011101110;
20'b01000001100110111111: color_data = 12'b111011101110;
20'b01000001100111000000: color_data = 12'b111011101110;
20'b01000001100111000001: color_data = 12'b111011101110;
20'b01000001100111000010: color_data = 12'b111011101110;
20'b01000001100111000011: color_data = 12'b111011101110;
20'b01000001100111000100: color_data = 12'b111011101110;
20'b01000001100111000101: color_data = 12'b111011101110;
20'b01000001100111000110: color_data = 12'b111011101110;
20'b01000001100111001000: color_data = 12'b111011101110;
20'b01000001100111001001: color_data = 12'b111011101110;
20'b01000001100111001010: color_data = 12'b111011101110;
20'b01000001100111001011: color_data = 12'b111011101110;
20'b01000001100111001100: color_data = 12'b111011101110;
20'b01000001100111001101: color_data = 12'b111011101110;
20'b01000001100111001110: color_data = 12'b111011101110;
20'b01000001100111001111: color_data = 12'b111011101110;
20'b01000001100111010000: color_data = 12'b111011101110;
20'b01000001100111010001: color_data = 12'b111011101110;
20'b01000001110010110111: color_data = 12'b111011101110;
20'b01000001110010111000: color_data = 12'b111011101110;
20'b01000001110010111001: color_data = 12'b111011101110;
20'b01000001110010111010: color_data = 12'b111011101110;
20'b01000001110010111011: color_data = 12'b111011101110;
20'b01000001110010111100: color_data = 12'b111011101110;
20'b01000001110010111101: color_data = 12'b111011101110;
20'b01000001110010111110: color_data = 12'b111011101110;
20'b01000001110010111111: color_data = 12'b111011101110;
20'b01000001110011000000: color_data = 12'b111011101110;
20'b01000001110011000010: color_data = 12'b111011101110;
20'b01000001110011000011: color_data = 12'b111011101110;
20'b01000001110011000100: color_data = 12'b111011101110;
20'b01000001110011000101: color_data = 12'b111011101110;
20'b01000001110011000110: color_data = 12'b111011101110;
20'b01000001110011000111: color_data = 12'b111011101110;
20'b01000001110011001000: color_data = 12'b111011101110;
20'b01000001110011001001: color_data = 12'b111011101110;
20'b01000001110011001010: color_data = 12'b111011101110;
20'b01000001110011001011: color_data = 12'b111011101110;
20'b01000001110011001101: color_data = 12'b111011101110;
20'b01000001110011001110: color_data = 12'b111011101110;
20'b01000001110011001111: color_data = 12'b111011101110;
20'b01000001110011010000: color_data = 12'b111011101110;
20'b01000001110011010001: color_data = 12'b111011101110;
20'b01000001110011010010: color_data = 12'b111011101110;
20'b01000001110011010011: color_data = 12'b111011101110;
20'b01000001110011010100: color_data = 12'b111011101110;
20'b01000001110011010101: color_data = 12'b111011101110;
20'b01000001110011010110: color_data = 12'b111011101110;
20'b01000001110011111000: color_data = 12'b000001111111;
20'b01000001110011111001: color_data = 12'b000001111111;
20'b01000001110011111010: color_data = 12'b000001111111;
20'b01000001110011111011: color_data = 12'b000001111111;
20'b01000001110011111100: color_data = 12'b000001111111;
20'b01000001110011111101: color_data = 12'b000001111111;
20'b01000001110011111110: color_data = 12'b000001111111;
20'b01000001110011111111: color_data = 12'b000001111111;
20'b01000001110100000000: color_data = 12'b000001111111;
20'b01000001110100000001: color_data = 12'b000001111111;
20'b01000001110101000100: color_data = 12'b000011110111;
20'b01000001110101000101: color_data = 12'b000011110111;
20'b01000001110101000110: color_data = 12'b000011110111;
20'b01000001110101000111: color_data = 12'b000011110111;
20'b01000001110101001000: color_data = 12'b000011110111;
20'b01000001110101001001: color_data = 12'b000011110111;
20'b01000001110101001010: color_data = 12'b000011110111;
20'b01000001110101001011: color_data = 12'b000011110111;
20'b01000001110101001100: color_data = 12'b000011110111;
20'b01000001110101001101: color_data = 12'b000011110111;
20'b01000001110101100101: color_data = 12'b111011101110;
20'b01000001110101100110: color_data = 12'b111011101110;
20'b01000001110101100111: color_data = 12'b111011101110;
20'b01000001110101101000: color_data = 12'b111011101110;
20'b01000001110101101001: color_data = 12'b111011101110;
20'b01000001110101101010: color_data = 12'b111011101110;
20'b01000001110101101011: color_data = 12'b111011101110;
20'b01000001110101101100: color_data = 12'b111011101110;
20'b01000001110101101101: color_data = 12'b111011101110;
20'b01000001110101101110: color_data = 12'b111011101110;
20'b01000001110101110000: color_data = 12'b111011101110;
20'b01000001110101110001: color_data = 12'b111011101110;
20'b01000001110101110010: color_data = 12'b111011101110;
20'b01000001110101110011: color_data = 12'b111011101110;
20'b01000001110101110100: color_data = 12'b111011101110;
20'b01000001110101110101: color_data = 12'b111011101110;
20'b01000001110101110110: color_data = 12'b111011101110;
20'b01000001110101110111: color_data = 12'b111011101110;
20'b01000001110101111000: color_data = 12'b111011101110;
20'b01000001110101111001: color_data = 12'b111011101110;
20'b01000001110101111011: color_data = 12'b111011101110;
20'b01000001110101111100: color_data = 12'b111011101110;
20'b01000001110101111101: color_data = 12'b111011101110;
20'b01000001110101111110: color_data = 12'b111011101110;
20'b01000001110101111111: color_data = 12'b111011101110;
20'b01000001110110000000: color_data = 12'b111011101110;
20'b01000001110110000001: color_data = 12'b111011101110;
20'b01000001110110000010: color_data = 12'b111011101110;
20'b01000001110110000011: color_data = 12'b111011101110;
20'b01000001110110000100: color_data = 12'b111011101110;
20'b01000001110110000110: color_data = 12'b111011101110;
20'b01000001110110000111: color_data = 12'b111011101110;
20'b01000001110110001000: color_data = 12'b111011101110;
20'b01000001110110001001: color_data = 12'b111011101110;
20'b01000001110110001010: color_data = 12'b111011101110;
20'b01000001110110001011: color_data = 12'b111011101110;
20'b01000001110110001100: color_data = 12'b111011101110;
20'b01000001110110001101: color_data = 12'b111011101110;
20'b01000001110110001110: color_data = 12'b111011101110;
20'b01000001110110001111: color_data = 12'b111011101110;
20'b01000001110110100111: color_data = 12'b111011101110;
20'b01000001110110101000: color_data = 12'b111011101110;
20'b01000001110110101001: color_data = 12'b111011101110;
20'b01000001110110101010: color_data = 12'b111011101110;
20'b01000001110110101011: color_data = 12'b111011101110;
20'b01000001110110101100: color_data = 12'b111011101110;
20'b01000001110110101101: color_data = 12'b111011101110;
20'b01000001110110101110: color_data = 12'b111011101110;
20'b01000001110110101111: color_data = 12'b111011101110;
20'b01000001110110110000: color_data = 12'b111011101110;
20'b01000001110110110010: color_data = 12'b111011101110;
20'b01000001110110110011: color_data = 12'b111011101110;
20'b01000001110110110100: color_data = 12'b111011101110;
20'b01000001110110110101: color_data = 12'b111011101110;
20'b01000001110110110110: color_data = 12'b111011101110;
20'b01000001110110110111: color_data = 12'b111011101110;
20'b01000001110110111000: color_data = 12'b111011101110;
20'b01000001110110111001: color_data = 12'b111011101110;
20'b01000001110110111010: color_data = 12'b111011101110;
20'b01000001110110111011: color_data = 12'b111011101110;
20'b01000001110110111101: color_data = 12'b111011101110;
20'b01000001110110111110: color_data = 12'b111011101110;
20'b01000001110110111111: color_data = 12'b111011101110;
20'b01000001110111000000: color_data = 12'b111011101110;
20'b01000001110111000001: color_data = 12'b111011101110;
20'b01000001110111000010: color_data = 12'b111011101110;
20'b01000001110111000011: color_data = 12'b111011101110;
20'b01000001110111000100: color_data = 12'b111011101110;
20'b01000001110111000101: color_data = 12'b111011101110;
20'b01000001110111000110: color_data = 12'b111011101110;
20'b01000001110111001000: color_data = 12'b111011101110;
20'b01000001110111001001: color_data = 12'b111011101110;
20'b01000001110111001010: color_data = 12'b111011101110;
20'b01000001110111001011: color_data = 12'b111011101110;
20'b01000001110111001100: color_data = 12'b111011101110;
20'b01000001110111001101: color_data = 12'b111011101110;
20'b01000001110111001110: color_data = 12'b111011101110;
20'b01000001110111001111: color_data = 12'b111011101110;
20'b01000001110111010000: color_data = 12'b111011101110;
20'b01000001110111010001: color_data = 12'b111011101110;
20'b01000010000010110111: color_data = 12'b111011101110;
20'b01000010000010111000: color_data = 12'b111011101110;
20'b01000010000010111001: color_data = 12'b111011101110;
20'b01000010000010111010: color_data = 12'b111011101110;
20'b01000010000010111011: color_data = 12'b111011101110;
20'b01000010000010111100: color_data = 12'b111011101110;
20'b01000010000010111101: color_data = 12'b111011101110;
20'b01000010000010111110: color_data = 12'b111011101110;
20'b01000010000010111111: color_data = 12'b111011101110;
20'b01000010000011000000: color_data = 12'b111011101110;
20'b01000010000011000010: color_data = 12'b111011101110;
20'b01000010000011000011: color_data = 12'b111011101110;
20'b01000010000011000100: color_data = 12'b111011101110;
20'b01000010000011000101: color_data = 12'b111011101110;
20'b01000010000011000110: color_data = 12'b111011101110;
20'b01000010000011000111: color_data = 12'b111011101110;
20'b01000010000011001000: color_data = 12'b111011101110;
20'b01000010000011001001: color_data = 12'b111011101110;
20'b01000010000011001010: color_data = 12'b111011101110;
20'b01000010000011001011: color_data = 12'b111011101110;
20'b01000010000011001101: color_data = 12'b111011101110;
20'b01000010000011001110: color_data = 12'b111011101110;
20'b01000010000011001111: color_data = 12'b111011101110;
20'b01000010000011010000: color_data = 12'b111011101110;
20'b01000010000011010001: color_data = 12'b111011101110;
20'b01000010000011010010: color_data = 12'b111011101110;
20'b01000010000011010011: color_data = 12'b111011101110;
20'b01000010000011010100: color_data = 12'b111011101110;
20'b01000010000011010101: color_data = 12'b111011101110;
20'b01000010000011010110: color_data = 12'b111011101110;
20'b01000010000011111000: color_data = 12'b000001111111;
20'b01000010000011111001: color_data = 12'b000001111111;
20'b01000010000011111010: color_data = 12'b000001111111;
20'b01000010000011111011: color_data = 12'b000001111111;
20'b01000010000011111100: color_data = 12'b000001111111;
20'b01000010000011111101: color_data = 12'b000001111111;
20'b01000010000011111110: color_data = 12'b000001111111;
20'b01000010000011111111: color_data = 12'b000001111111;
20'b01000010000100000000: color_data = 12'b000001111111;
20'b01000010000100000001: color_data = 12'b000001111111;
20'b01000010000101000100: color_data = 12'b000011110111;
20'b01000010000101000101: color_data = 12'b000011110111;
20'b01000010000101000110: color_data = 12'b000011110111;
20'b01000010000101000111: color_data = 12'b000011110111;
20'b01000010000101001000: color_data = 12'b000011110111;
20'b01000010000101001001: color_data = 12'b000011110111;
20'b01000010000101001010: color_data = 12'b000011110111;
20'b01000010000101001011: color_data = 12'b000011110111;
20'b01000010000101001100: color_data = 12'b000011110111;
20'b01000010000101001101: color_data = 12'b000011110111;
20'b01000010000101100101: color_data = 12'b111011101110;
20'b01000010000101100110: color_data = 12'b111011101110;
20'b01000010000101100111: color_data = 12'b111011101110;
20'b01000010000101101000: color_data = 12'b111011101110;
20'b01000010000101101001: color_data = 12'b111011101110;
20'b01000010000101101010: color_data = 12'b111011101110;
20'b01000010000101101011: color_data = 12'b111011101110;
20'b01000010000101101100: color_data = 12'b111011101110;
20'b01000010000101101101: color_data = 12'b111011101110;
20'b01000010000101101110: color_data = 12'b111011101110;
20'b01000010000101110000: color_data = 12'b111011101110;
20'b01000010000101110001: color_data = 12'b111011101110;
20'b01000010000101110010: color_data = 12'b111011101110;
20'b01000010000101110011: color_data = 12'b111011101110;
20'b01000010000101110100: color_data = 12'b111011101110;
20'b01000010000101110101: color_data = 12'b111011101110;
20'b01000010000101110110: color_data = 12'b111011101110;
20'b01000010000101110111: color_data = 12'b111011101110;
20'b01000010000101111000: color_data = 12'b111011101110;
20'b01000010000101111001: color_data = 12'b111011101110;
20'b01000010000101111011: color_data = 12'b111011101110;
20'b01000010000101111100: color_data = 12'b111011101110;
20'b01000010000101111101: color_data = 12'b111011101110;
20'b01000010000101111110: color_data = 12'b111011101110;
20'b01000010000101111111: color_data = 12'b111011101110;
20'b01000010000110000000: color_data = 12'b111011101110;
20'b01000010000110000001: color_data = 12'b111011101110;
20'b01000010000110000010: color_data = 12'b111011101110;
20'b01000010000110000011: color_data = 12'b111011101110;
20'b01000010000110000100: color_data = 12'b111011101110;
20'b01000010000110000110: color_data = 12'b111011101110;
20'b01000010000110000111: color_data = 12'b111011101110;
20'b01000010000110001000: color_data = 12'b111011101110;
20'b01000010000110001001: color_data = 12'b111011101110;
20'b01000010000110001010: color_data = 12'b111011101110;
20'b01000010000110001011: color_data = 12'b111011101110;
20'b01000010000110001100: color_data = 12'b111011101110;
20'b01000010000110001101: color_data = 12'b111011101110;
20'b01000010000110001110: color_data = 12'b111011101110;
20'b01000010000110001111: color_data = 12'b111011101110;
20'b01000010000110100111: color_data = 12'b111011101110;
20'b01000010000110101000: color_data = 12'b111011101110;
20'b01000010000110101001: color_data = 12'b111011101110;
20'b01000010000110101010: color_data = 12'b111011101110;
20'b01000010000110101011: color_data = 12'b111011101110;
20'b01000010000110101100: color_data = 12'b111011101110;
20'b01000010000110101101: color_data = 12'b111011101110;
20'b01000010000110101110: color_data = 12'b111011101110;
20'b01000010000110101111: color_data = 12'b111011101110;
20'b01000010000110110000: color_data = 12'b111011101110;
20'b01000010000110110010: color_data = 12'b111011101110;
20'b01000010000110110011: color_data = 12'b111011101110;
20'b01000010000110110100: color_data = 12'b111011101110;
20'b01000010000110110101: color_data = 12'b111011101110;
20'b01000010000110110110: color_data = 12'b111011101110;
20'b01000010000110110111: color_data = 12'b111011101110;
20'b01000010000110111000: color_data = 12'b111011101110;
20'b01000010000110111001: color_data = 12'b111011101110;
20'b01000010000110111010: color_data = 12'b111011101110;
20'b01000010000110111011: color_data = 12'b111011101110;
20'b01000010000110111101: color_data = 12'b111011101110;
20'b01000010000110111110: color_data = 12'b111011101110;
20'b01000010000110111111: color_data = 12'b111011101110;
20'b01000010000111000000: color_data = 12'b111011101110;
20'b01000010000111000001: color_data = 12'b111011101110;
20'b01000010000111000010: color_data = 12'b111011101110;
20'b01000010000111000011: color_data = 12'b111011101110;
20'b01000010000111000100: color_data = 12'b111011101110;
20'b01000010000111000101: color_data = 12'b111011101110;
20'b01000010000111000110: color_data = 12'b111011101110;
20'b01000010000111001000: color_data = 12'b111011101110;
20'b01000010000111001001: color_data = 12'b111011101110;
20'b01000010000111001010: color_data = 12'b111011101110;
20'b01000010000111001011: color_data = 12'b111011101110;
20'b01000010000111001100: color_data = 12'b111011101110;
20'b01000010000111001101: color_data = 12'b111011101110;
20'b01000010000111001110: color_data = 12'b111011101110;
20'b01000010000111001111: color_data = 12'b111011101110;
20'b01000010000111010000: color_data = 12'b111011101110;
20'b01000010000111010001: color_data = 12'b111011101110;
20'b01000010010010110111: color_data = 12'b111011101110;
20'b01000010010010111000: color_data = 12'b111011101110;
20'b01000010010010111001: color_data = 12'b111011101110;
20'b01000010010010111010: color_data = 12'b111011101110;
20'b01000010010010111011: color_data = 12'b111011101110;
20'b01000010010010111100: color_data = 12'b111011101110;
20'b01000010010010111101: color_data = 12'b111011101110;
20'b01000010010010111110: color_data = 12'b111011101110;
20'b01000010010010111111: color_data = 12'b111011101110;
20'b01000010010011000000: color_data = 12'b111011101110;
20'b01000010010011000010: color_data = 12'b111011101110;
20'b01000010010011000011: color_data = 12'b111011101110;
20'b01000010010011000100: color_data = 12'b111011101110;
20'b01000010010011000101: color_data = 12'b111011101110;
20'b01000010010011000110: color_data = 12'b111011101110;
20'b01000010010011000111: color_data = 12'b111011101110;
20'b01000010010011001000: color_data = 12'b111011101110;
20'b01000010010011001001: color_data = 12'b111011101110;
20'b01000010010011001010: color_data = 12'b111011101110;
20'b01000010010011001011: color_data = 12'b111011101110;
20'b01000010010011001101: color_data = 12'b111011101110;
20'b01000010010011001110: color_data = 12'b111011101110;
20'b01000010010011001111: color_data = 12'b111011101110;
20'b01000010010011010000: color_data = 12'b111011101110;
20'b01000010010011010001: color_data = 12'b111011101110;
20'b01000010010011010010: color_data = 12'b111011101110;
20'b01000010010011010011: color_data = 12'b111011101110;
20'b01000010010011010100: color_data = 12'b111011101110;
20'b01000010010011010101: color_data = 12'b111011101110;
20'b01000010010011010110: color_data = 12'b111011101110;
20'b01000010010011111000: color_data = 12'b000001111111;
20'b01000010010011111001: color_data = 12'b000001111111;
20'b01000010010011111010: color_data = 12'b000001111111;
20'b01000010010011111011: color_data = 12'b000001111111;
20'b01000010010011111100: color_data = 12'b000001111111;
20'b01000010010011111101: color_data = 12'b000001111111;
20'b01000010010011111110: color_data = 12'b000001111111;
20'b01000010010011111111: color_data = 12'b000001111111;
20'b01000010010100000000: color_data = 12'b000001111111;
20'b01000010010100000001: color_data = 12'b000001111111;
20'b01000010010101000100: color_data = 12'b000011110111;
20'b01000010010101000101: color_data = 12'b000011110111;
20'b01000010010101000110: color_data = 12'b000011110111;
20'b01000010010101000111: color_data = 12'b000011110111;
20'b01000010010101001000: color_data = 12'b000011110111;
20'b01000010010101001001: color_data = 12'b000011110111;
20'b01000010010101001010: color_data = 12'b000011110111;
20'b01000010010101001011: color_data = 12'b000011110111;
20'b01000010010101001100: color_data = 12'b000011110111;
20'b01000010010101001101: color_data = 12'b000011110111;
20'b01000010010101100101: color_data = 12'b111011101110;
20'b01000010010101100110: color_data = 12'b111011101110;
20'b01000010010101100111: color_data = 12'b111011101110;
20'b01000010010101101000: color_data = 12'b111011101110;
20'b01000010010101101001: color_data = 12'b111011101110;
20'b01000010010101101010: color_data = 12'b111011101110;
20'b01000010010101101011: color_data = 12'b111011101110;
20'b01000010010101101100: color_data = 12'b111011101110;
20'b01000010010101101101: color_data = 12'b111011101110;
20'b01000010010101101110: color_data = 12'b111011101110;
20'b01000010010101110000: color_data = 12'b111011101110;
20'b01000010010101110001: color_data = 12'b111011101110;
20'b01000010010101110010: color_data = 12'b111011101110;
20'b01000010010101110011: color_data = 12'b111011101110;
20'b01000010010101110100: color_data = 12'b111011101110;
20'b01000010010101110101: color_data = 12'b111011101110;
20'b01000010010101110110: color_data = 12'b111011101110;
20'b01000010010101110111: color_data = 12'b111011101110;
20'b01000010010101111000: color_data = 12'b111011101110;
20'b01000010010101111001: color_data = 12'b111011101110;
20'b01000010010101111011: color_data = 12'b111011101110;
20'b01000010010101111100: color_data = 12'b111011101110;
20'b01000010010101111101: color_data = 12'b111011101110;
20'b01000010010101111110: color_data = 12'b111011101110;
20'b01000010010101111111: color_data = 12'b111011101110;
20'b01000010010110000000: color_data = 12'b111011101110;
20'b01000010010110000001: color_data = 12'b111011101110;
20'b01000010010110000010: color_data = 12'b111011101110;
20'b01000010010110000011: color_data = 12'b111011101110;
20'b01000010010110000100: color_data = 12'b111011101110;
20'b01000010010110000110: color_data = 12'b111011101110;
20'b01000010010110000111: color_data = 12'b111011101110;
20'b01000010010110001000: color_data = 12'b111011101110;
20'b01000010010110001001: color_data = 12'b111011101110;
20'b01000010010110001010: color_data = 12'b111011101110;
20'b01000010010110001011: color_data = 12'b111011101110;
20'b01000010010110001100: color_data = 12'b111011101110;
20'b01000010010110001101: color_data = 12'b111011101110;
20'b01000010010110001110: color_data = 12'b111011101110;
20'b01000010010110001111: color_data = 12'b111011101110;
20'b01000010010110100111: color_data = 12'b111011101110;
20'b01000010010110101000: color_data = 12'b111011101110;
20'b01000010010110101001: color_data = 12'b111011101110;
20'b01000010010110101010: color_data = 12'b111011101110;
20'b01000010010110101011: color_data = 12'b111011101110;
20'b01000010010110101100: color_data = 12'b111011101110;
20'b01000010010110101101: color_data = 12'b111011101110;
20'b01000010010110101110: color_data = 12'b111011101110;
20'b01000010010110101111: color_data = 12'b111011101110;
20'b01000010010110110000: color_data = 12'b111011101110;
20'b01000010010110110010: color_data = 12'b111011101110;
20'b01000010010110110011: color_data = 12'b111011101110;
20'b01000010010110110100: color_data = 12'b111011101110;
20'b01000010010110110101: color_data = 12'b111011101110;
20'b01000010010110110110: color_data = 12'b111011101110;
20'b01000010010110110111: color_data = 12'b111011101110;
20'b01000010010110111000: color_data = 12'b111011101110;
20'b01000010010110111001: color_data = 12'b111011101110;
20'b01000010010110111010: color_data = 12'b111011101110;
20'b01000010010110111011: color_data = 12'b111011101110;
20'b01000010010110111101: color_data = 12'b111011101110;
20'b01000010010110111110: color_data = 12'b111011101110;
20'b01000010010110111111: color_data = 12'b111011101110;
20'b01000010010111000000: color_data = 12'b111011101110;
20'b01000010010111000001: color_data = 12'b111011101110;
20'b01000010010111000010: color_data = 12'b111011101110;
20'b01000010010111000011: color_data = 12'b111011101110;
20'b01000010010111000100: color_data = 12'b111011101110;
20'b01000010010111000101: color_data = 12'b111011101110;
20'b01000010010111000110: color_data = 12'b111011101110;
20'b01000010010111001000: color_data = 12'b111011101110;
20'b01000010010111001001: color_data = 12'b111011101110;
20'b01000010010111001010: color_data = 12'b111011101110;
20'b01000010010111001011: color_data = 12'b111011101110;
20'b01000010010111001100: color_data = 12'b111011101110;
20'b01000010010111001101: color_data = 12'b111011101110;
20'b01000010010111001110: color_data = 12'b111011101110;
20'b01000010010111001111: color_data = 12'b111011101110;
20'b01000010010111010000: color_data = 12'b111011101110;
20'b01000010010111010001: color_data = 12'b111011101110;
20'b01000010110010010110: color_data = 12'b111011101110;
20'b01000010110010010111: color_data = 12'b111011101110;
20'b01000010110010011000: color_data = 12'b111011101110;
20'b01000010110010011001: color_data = 12'b111011101110;
20'b01000010110010011010: color_data = 12'b111011101110;
20'b01000010110010011011: color_data = 12'b111011101110;
20'b01000010110010011100: color_data = 12'b111011101110;
20'b01000010110010011101: color_data = 12'b111011101110;
20'b01000010110010011110: color_data = 12'b111011101110;
20'b01000010110010011111: color_data = 12'b111011101110;
20'b01000010110011001101: color_data = 12'b111011101110;
20'b01000010110011001110: color_data = 12'b111011101110;
20'b01000010110011001111: color_data = 12'b111011101110;
20'b01000010110011010000: color_data = 12'b111011101110;
20'b01000010110011010001: color_data = 12'b111011101110;
20'b01000010110011010010: color_data = 12'b111011101110;
20'b01000010110011010011: color_data = 12'b111011101110;
20'b01000010110011010100: color_data = 12'b111011101110;
20'b01000010110011010101: color_data = 12'b111011101110;
20'b01000010110011010110: color_data = 12'b111011101110;
20'b01000010110011011000: color_data = 12'b111011101110;
20'b01000010110011011001: color_data = 12'b111011101110;
20'b01000010110011011010: color_data = 12'b111011101110;
20'b01000010110011011011: color_data = 12'b111011101110;
20'b01000010110011011100: color_data = 12'b111011101110;
20'b01000010110011011101: color_data = 12'b111011101110;
20'b01000010110011011110: color_data = 12'b111011101110;
20'b01000010110011011111: color_data = 12'b111011101110;
20'b01000010110011100000: color_data = 12'b111011101110;
20'b01000010110011100001: color_data = 12'b111011101110;
20'b01000010110011101101: color_data = 12'b111011101110;
20'b01000010110011101110: color_data = 12'b111011101110;
20'b01000010110011101111: color_data = 12'b111011101110;
20'b01000010110011110000: color_data = 12'b111011101110;
20'b01000010110011110001: color_data = 12'b111011101110;
20'b01000010110011110010: color_data = 12'b111011101110;
20'b01000010110011110011: color_data = 12'b111011101110;
20'b01000010110011110100: color_data = 12'b111011101110;
20'b01000010110011110101: color_data = 12'b111011101110;
20'b01000010110011110110: color_data = 12'b111011101110;
20'b01000010110101001111: color_data = 12'b111011101110;
20'b01000010110101010000: color_data = 12'b111011101110;
20'b01000010110101010001: color_data = 12'b111011101110;
20'b01000010110101010010: color_data = 12'b111011101110;
20'b01000010110101010011: color_data = 12'b111011101110;
20'b01000010110101010100: color_data = 12'b111011101110;
20'b01000010110101010101: color_data = 12'b111011101110;
20'b01000010110101010110: color_data = 12'b111011101110;
20'b01000010110101010111: color_data = 12'b111011101110;
20'b01000010110101011000: color_data = 12'b111011101110;
20'b01000010110110011100: color_data = 12'b111011101110;
20'b01000010110110011101: color_data = 12'b111011101110;
20'b01000010110110011110: color_data = 12'b111011101110;
20'b01000010110110011111: color_data = 12'b111011101110;
20'b01000010110110100000: color_data = 12'b111011101110;
20'b01000010110110100001: color_data = 12'b111011101110;
20'b01000010110110100010: color_data = 12'b111011101110;
20'b01000010110110100011: color_data = 12'b111011101110;
20'b01000010110110100100: color_data = 12'b111011101110;
20'b01000010110110100101: color_data = 12'b111011101110;
20'b01000010110110100111: color_data = 12'b111011101110;
20'b01000010110110101000: color_data = 12'b111011101110;
20'b01000010110110101001: color_data = 12'b111011101110;
20'b01000010110110101010: color_data = 12'b111011101110;
20'b01000010110110101011: color_data = 12'b111011101110;
20'b01000010110110101100: color_data = 12'b111011101110;
20'b01000010110110101101: color_data = 12'b111011101110;
20'b01000010110110101110: color_data = 12'b111011101110;
20'b01000010110110101111: color_data = 12'b111011101110;
20'b01000010110110110000: color_data = 12'b111011101110;
20'b01000011000010010110: color_data = 12'b111011101110;
20'b01000011000010010111: color_data = 12'b111011101110;
20'b01000011000010011000: color_data = 12'b111011101110;
20'b01000011000010011001: color_data = 12'b111011101110;
20'b01000011000010011010: color_data = 12'b111011101110;
20'b01000011000010011011: color_data = 12'b111011101110;
20'b01000011000010011100: color_data = 12'b111011101110;
20'b01000011000010011101: color_data = 12'b111011101110;
20'b01000011000010011110: color_data = 12'b111011101110;
20'b01000011000010011111: color_data = 12'b111011101110;
20'b01000011000011001101: color_data = 12'b111011101110;
20'b01000011000011001110: color_data = 12'b111011101110;
20'b01000011000011001111: color_data = 12'b111011101110;
20'b01000011000011010000: color_data = 12'b111011101110;
20'b01000011000011010001: color_data = 12'b111011101110;
20'b01000011000011010010: color_data = 12'b111011101110;
20'b01000011000011010011: color_data = 12'b111011101110;
20'b01000011000011010100: color_data = 12'b111011101110;
20'b01000011000011010101: color_data = 12'b111011101110;
20'b01000011000011010110: color_data = 12'b111011101110;
20'b01000011000011011000: color_data = 12'b111011101110;
20'b01000011000011011001: color_data = 12'b111011101110;
20'b01000011000011011010: color_data = 12'b111011101110;
20'b01000011000011011011: color_data = 12'b111011101110;
20'b01000011000011011100: color_data = 12'b111011101110;
20'b01000011000011011101: color_data = 12'b111011101110;
20'b01000011000011011110: color_data = 12'b111011101110;
20'b01000011000011011111: color_data = 12'b111011101110;
20'b01000011000011100000: color_data = 12'b111011101110;
20'b01000011000011100001: color_data = 12'b111011101110;
20'b01000011000011101101: color_data = 12'b111011101110;
20'b01000011000011101110: color_data = 12'b111011101110;
20'b01000011000011101111: color_data = 12'b111011101110;
20'b01000011000011110000: color_data = 12'b111011101110;
20'b01000011000011110001: color_data = 12'b111011101110;
20'b01000011000011110010: color_data = 12'b111011101110;
20'b01000011000011110011: color_data = 12'b111011101110;
20'b01000011000011110100: color_data = 12'b111011101110;
20'b01000011000011110101: color_data = 12'b111011101110;
20'b01000011000011110110: color_data = 12'b111011101110;
20'b01000011000101001111: color_data = 12'b111011101110;
20'b01000011000101010000: color_data = 12'b111011101110;
20'b01000011000101010001: color_data = 12'b111011101110;
20'b01000011000101010010: color_data = 12'b111011101110;
20'b01000011000101010011: color_data = 12'b111011101110;
20'b01000011000101010100: color_data = 12'b111011101110;
20'b01000011000101010101: color_data = 12'b111011101110;
20'b01000011000101010110: color_data = 12'b111011101110;
20'b01000011000101010111: color_data = 12'b111011101110;
20'b01000011000101011000: color_data = 12'b111011101110;
20'b01000011000110011100: color_data = 12'b111011101110;
20'b01000011000110011101: color_data = 12'b111011101110;
20'b01000011000110011110: color_data = 12'b111011101110;
20'b01000011000110011111: color_data = 12'b111011101110;
20'b01000011000110100000: color_data = 12'b111011101110;
20'b01000011000110100001: color_data = 12'b111011101110;
20'b01000011000110100010: color_data = 12'b111011101110;
20'b01000011000110100011: color_data = 12'b111011101110;
20'b01000011000110100100: color_data = 12'b111011101110;
20'b01000011000110100101: color_data = 12'b111011101110;
20'b01000011000110100111: color_data = 12'b111011101110;
20'b01000011000110101000: color_data = 12'b111011101110;
20'b01000011000110101001: color_data = 12'b111011101110;
20'b01000011000110101010: color_data = 12'b111011101110;
20'b01000011000110101011: color_data = 12'b111011101110;
20'b01000011000110101100: color_data = 12'b111011101110;
20'b01000011000110101101: color_data = 12'b111011101110;
20'b01000011000110101110: color_data = 12'b111011101110;
20'b01000011000110101111: color_data = 12'b111011101110;
20'b01000011000110110000: color_data = 12'b111011101110;
20'b01000011010010010110: color_data = 12'b111011101110;
20'b01000011010010010111: color_data = 12'b111011101110;
20'b01000011010010011000: color_data = 12'b111011101110;
20'b01000011010010011001: color_data = 12'b111011101110;
20'b01000011010010011010: color_data = 12'b111011101110;
20'b01000011010010011011: color_data = 12'b111011101110;
20'b01000011010010011100: color_data = 12'b111011101110;
20'b01000011010010011101: color_data = 12'b111011101110;
20'b01000011010010011110: color_data = 12'b111011101110;
20'b01000011010010011111: color_data = 12'b111011101110;
20'b01000011010011001101: color_data = 12'b111011101110;
20'b01000011010011001110: color_data = 12'b111011101110;
20'b01000011010011001111: color_data = 12'b111011101110;
20'b01000011010011010000: color_data = 12'b111011101110;
20'b01000011010011010001: color_data = 12'b111011101110;
20'b01000011010011010010: color_data = 12'b111011101110;
20'b01000011010011010011: color_data = 12'b111011101110;
20'b01000011010011010100: color_data = 12'b111011101110;
20'b01000011010011010101: color_data = 12'b111011101110;
20'b01000011010011010110: color_data = 12'b111011101110;
20'b01000011010011011000: color_data = 12'b111011101110;
20'b01000011010011011001: color_data = 12'b111011101110;
20'b01000011010011011010: color_data = 12'b111011101110;
20'b01000011010011011011: color_data = 12'b111011101110;
20'b01000011010011011100: color_data = 12'b111011101110;
20'b01000011010011011101: color_data = 12'b111011101110;
20'b01000011010011011110: color_data = 12'b111011101110;
20'b01000011010011011111: color_data = 12'b111011101110;
20'b01000011010011100000: color_data = 12'b111011101110;
20'b01000011010011100001: color_data = 12'b111011101110;
20'b01000011010011101101: color_data = 12'b111011101110;
20'b01000011010011101110: color_data = 12'b111011101110;
20'b01000011010011101111: color_data = 12'b111011101110;
20'b01000011010011110000: color_data = 12'b111011101110;
20'b01000011010011110001: color_data = 12'b111011101110;
20'b01000011010011110010: color_data = 12'b111011101110;
20'b01000011010011110011: color_data = 12'b111011101110;
20'b01000011010011110100: color_data = 12'b111011101110;
20'b01000011010011110101: color_data = 12'b111011101110;
20'b01000011010011110110: color_data = 12'b111011101110;
20'b01000011010101001111: color_data = 12'b111011101110;
20'b01000011010101010000: color_data = 12'b111011101110;
20'b01000011010101010001: color_data = 12'b111011101110;
20'b01000011010101010010: color_data = 12'b111011101110;
20'b01000011010101010011: color_data = 12'b111011101110;
20'b01000011010101010100: color_data = 12'b111011101110;
20'b01000011010101010101: color_data = 12'b111011101110;
20'b01000011010101010110: color_data = 12'b111011101110;
20'b01000011010101010111: color_data = 12'b111011101110;
20'b01000011010101011000: color_data = 12'b111011101110;
20'b01000011010110011100: color_data = 12'b111011101110;
20'b01000011010110011101: color_data = 12'b111011101110;
20'b01000011010110011110: color_data = 12'b111011101110;
20'b01000011010110011111: color_data = 12'b111011101110;
20'b01000011010110100000: color_data = 12'b111011101110;
20'b01000011010110100001: color_data = 12'b111011101110;
20'b01000011010110100010: color_data = 12'b111011101110;
20'b01000011010110100011: color_data = 12'b111011101110;
20'b01000011010110100100: color_data = 12'b111011101110;
20'b01000011010110100101: color_data = 12'b111011101110;
20'b01000011010110100111: color_data = 12'b111011101110;
20'b01000011010110101000: color_data = 12'b111011101110;
20'b01000011010110101001: color_data = 12'b111011101110;
20'b01000011010110101010: color_data = 12'b111011101110;
20'b01000011010110101011: color_data = 12'b111011101110;
20'b01000011010110101100: color_data = 12'b111011101110;
20'b01000011010110101101: color_data = 12'b111011101110;
20'b01000011010110101110: color_data = 12'b111011101110;
20'b01000011010110101111: color_data = 12'b111011101110;
20'b01000011010110110000: color_data = 12'b111011101110;
20'b01000011100010010110: color_data = 12'b111011101110;
20'b01000011100010010111: color_data = 12'b111011101110;
20'b01000011100010011000: color_data = 12'b111011101110;
20'b01000011100010011001: color_data = 12'b111011101110;
20'b01000011100010011010: color_data = 12'b111011101110;
20'b01000011100010011011: color_data = 12'b111011101110;
20'b01000011100010011100: color_data = 12'b111011101110;
20'b01000011100010011101: color_data = 12'b111011101110;
20'b01000011100010011110: color_data = 12'b111011101110;
20'b01000011100010011111: color_data = 12'b111011101110;
20'b01000011100011001101: color_data = 12'b111011101110;
20'b01000011100011001110: color_data = 12'b111011101110;
20'b01000011100011001111: color_data = 12'b111011101110;
20'b01000011100011010000: color_data = 12'b111011101110;
20'b01000011100011010001: color_data = 12'b111011101110;
20'b01000011100011010010: color_data = 12'b111011101110;
20'b01000011100011010011: color_data = 12'b111011101110;
20'b01000011100011010100: color_data = 12'b111011101110;
20'b01000011100011010101: color_data = 12'b111011101110;
20'b01000011100011010110: color_data = 12'b111011101110;
20'b01000011100011011000: color_data = 12'b111011101110;
20'b01000011100011011001: color_data = 12'b111011101110;
20'b01000011100011011010: color_data = 12'b111011101110;
20'b01000011100011011011: color_data = 12'b111011101110;
20'b01000011100011011100: color_data = 12'b111011101110;
20'b01000011100011011101: color_data = 12'b111011101110;
20'b01000011100011011110: color_data = 12'b111011101110;
20'b01000011100011011111: color_data = 12'b111011101110;
20'b01000011100011100000: color_data = 12'b111011101110;
20'b01000011100011100001: color_data = 12'b111011101110;
20'b01000011100011101101: color_data = 12'b111011101110;
20'b01000011100011101110: color_data = 12'b111011101110;
20'b01000011100011101111: color_data = 12'b111011101110;
20'b01000011100011110000: color_data = 12'b111011101110;
20'b01000011100011110001: color_data = 12'b111011101110;
20'b01000011100011110010: color_data = 12'b111011101110;
20'b01000011100011110011: color_data = 12'b111011101110;
20'b01000011100011110100: color_data = 12'b111011101110;
20'b01000011100011110101: color_data = 12'b111011101110;
20'b01000011100011110110: color_data = 12'b111011101110;
20'b01000011100101001111: color_data = 12'b111011101110;
20'b01000011100101010000: color_data = 12'b111011101110;
20'b01000011100101010001: color_data = 12'b111011101110;
20'b01000011100101010010: color_data = 12'b111011101110;
20'b01000011100101010011: color_data = 12'b111011101110;
20'b01000011100101010100: color_data = 12'b111011101110;
20'b01000011100101010101: color_data = 12'b111011101110;
20'b01000011100101010110: color_data = 12'b111011101110;
20'b01000011100101010111: color_data = 12'b111011101110;
20'b01000011100101011000: color_data = 12'b111011101110;
20'b01000011100110011100: color_data = 12'b111011101110;
20'b01000011100110011101: color_data = 12'b111011101110;
20'b01000011100110011110: color_data = 12'b111011101110;
20'b01000011100110011111: color_data = 12'b111011101110;
20'b01000011100110100000: color_data = 12'b111011101110;
20'b01000011100110100001: color_data = 12'b111011101110;
20'b01000011100110100010: color_data = 12'b111011101110;
20'b01000011100110100011: color_data = 12'b111011101110;
20'b01000011100110100100: color_data = 12'b111011101110;
20'b01000011100110100101: color_data = 12'b111011101110;
20'b01000011100110100111: color_data = 12'b111011101110;
20'b01000011100110101000: color_data = 12'b111011101110;
20'b01000011100110101001: color_data = 12'b111011101110;
20'b01000011100110101010: color_data = 12'b111011101110;
20'b01000011100110101011: color_data = 12'b111011101110;
20'b01000011100110101100: color_data = 12'b111011101110;
20'b01000011100110101101: color_data = 12'b111011101110;
20'b01000011100110101110: color_data = 12'b111011101110;
20'b01000011100110101111: color_data = 12'b111011101110;
20'b01000011100110110000: color_data = 12'b111011101110;
20'b01000011110010010110: color_data = 12'b111011101110;
20'b01000011110010010111: color_data = 12'b111011101110;
20'b01000011110010011000: color_data = 12'b111011101110;
20'b01000011110010011001: color_data = 12'b111011101110;
20'b01000011110010011010: color_data = 12'b111011101110;
20'b01000011110010011011: color_data = 12'b111011101110;
20'b01000011110010011100: color_data = 12'b111011101110;
20'b01000011110010011101: color_data = 12'b111011101110;
20'b01000011110010011110: color_data = 12'b111011101110;
20'b01000011110010011111: color_data = 12'b111011101110;
20'b01000011110011001101: color_data = 12'b111011101110;
20'b01000011110011001110: color_data = 12'b111011101110;
20'b01000011110011001111: color_data = 12'b111011101110;
20'b01000011110011010000: color_data = 12'b111011101110;
20'b01000011110011010001: color_data = 12'b111011101110;
20'b01000011110011010010: color_data = 12'b111011101110;
20'b01000011110011010011: color_data = 12'b111011101110;
20'b01000011110011010100: color_data = 12'b111011101110;
20'b01000011110011010101: color_data = 12'b111011101110;
20'b01000011110011010110: color_data = 12'b111011101110;
20'b01000011110011011000: color_data = 12'b111011101110;
20'b01000011110011011001: color_data = 12'b111011101110;
20'b01000011110011011010: color_data = 12'b111011101110;
20'b01000011110011011011: color_data = 12'b111011101110;
20'b01000011110011011100: color_data = 12'b111011101110;
20'b01000011110011011101: color_data = 12'b111011101110;
20'b01000011110011011110: color_data = 12'b111011101110;
20'b01000011110011011111: color_data = 12'b111011101110;
20'b01000011110011100000: color_data = 12'b111011101110;
20'b01000011110011100001: color_data = 12'b111011101110;
20'b01000011110011101101: color_data = 12'b111011101110;
20'b01000011110011101110: color_data = 12'b111011101110;
20'b01000011110011101111: color_data = 12'b111011101110;
20'b01000011110011110000: color_data = 12'b111011101110;
20'b01000011110011110001: color_data = 12'b111011101110;
20'b01000011110011110010: color_data = 12'b111011101110;
20'b01000011110011110011: color_data = 12'b111011101110;
20'b01000011110011110100: color_data = 12'b111011101110;
20'b01000011110011110101: color_data = 12'b111011101110;
20'b01000011110011110110: color_data = 12'b111011101110;
20'b01000011110101001111: color_data = 12'b111011101110;
20'b01000011110101010000: color_data = 12'b111011101110;
20'b01000011110101010001: color_data = 12'b111011101110;
20'b01000011110101010010: color_data = 12'b111011101110;
20'b01000011110101010011: color_data = 12'b111011101110;
20'b01000011110101010100: color_data = 12'b111011101110;
20'b01000011110101010101: color_data = 12'b111011101110;
20'b01000011110101010110: color_data = 12'b111011101110;
20'b01000011110101010111: color_data = 12'b111011101110;
20'b01000011110101011000: color_data = 12'b111011101110;
20'b01000011110110011100: color_data = 12'b111011101110;
20'b01000011110110011101: color_data = 12'b111011101110;
20'b01000011110110011110: color_data = 12'b111011101110;
20'b01000011110110011111: color_data = 12'b111011101110;
20'b01000011110110100000: color_data = 12'b111011101110;
20'b01000011110110100001: color_data = 12'b111011101110;
20'b01000011110110100010: color_data = 12'b111011101110;
20'b01000011110110100011: color_data = 12'b111011101110;
20'b01000011110110100100: color_data = 12'b111011101110;
20'b01000011110110100101: color_data = 12'b111011101110;
20'b01000011110110100111: color_data = 12'b111011101110;
20'b01000011110110101000: color_data = 12'b111011101110;
20'b01000011110110101001: color_data = 12'b111011101110;
20'b01000011110110101010: color_data = 12'b111011101110;
20'b01000011110110101011: color_data = 12'b111011101110;
20'b01000011110110101100: color_data = 12'b111011101110;
20'b01000011110110101101: color_data = 12'b111011101110;
20'b01000011110110101110: color_data = 12'b111011101110;
20'b01000011110110101111: color_data = 12'b111011101110;
20'b01000011110110110000: color_data = 12'b111011101110;
20'b01000100000010010110: color_data = 12'b111011101110;
20'b01000100000010010111: color_data = 12'b111011101110;
20'b01000100000010011000: color_data = 12'b111011101110;
20'b01000100000010011001: color_data = 12'b111011101110;
20'b01000100000010011010: color_data = 12'b111011101110;
20'b01000100000010011011: color_data = 12'b111011101110;
20'b01000100000010011100: color_data = 12'b111011101110;
20'b01000100000010011101: color_data = 12'b111011101110;
20'b01000100000010011110: color_data = 12'b111011101110;
20'b01000100000010011111: color_data = 12'b111011101110;
20'b01000100000011001101: color_data = 12'b111011101110;
20'b01000100000011001110: color_data = 12'b111011101110;
20'b01000100000011001111: color_data = 12'b111011101110;
20'b01000100000011010000: color_data = 12'b111011101110;
20'b01000100000011010001: color_data = 12'b111011101110;
20'b01000100000011010010: color_data = 12'b111011101110;
20'b01000100000011010011: color_data = 12'b111011101110;
20'b01000100000011010100: color_data = 12'b111011101110;
20'b01000100000011010101: color_data = 12'b111011101110;
20'b01000100000011010110: color_data = 12'b111011101110;
20'b01000100000011011000: color_data = 12'b111011101110;
20'b01000100000011011001: color_data = 12'b111011101110;
20'b01000100000011011010: color_data = 12'b111011101110;
20'b01000100000011011011: color_data = 12'b111011101110;
20'b01000100000011011100: color_data = 12'b111011101110;
20'b01000100000011011101: color_data = 12'b111011101110;
20'b01000100000011011110: color_data = 12'b111011101110;
20'b01000100000011011111: color_data = 12'b111011101110;
20'b01000100000011100000: color_data = 12'b111011101110;
20'b01000100000011100001: color_data = 12'b111011101110;
20'b01000100000011101101: color_data = 12'b111011101110;
20'b01000100000011101110: color_data = 12'b111011101110;
20'b01000100000011101111: color_data = 12'b111011101110;
20'b01000100000011110000: color_data = 12'b111011101110;
20'b01000100000011110001: color_data = 12'b111011101110;
20'b01000100000011110010: color_data = 12'b111011101110;
20'b01000100000011110011: color_data = 12'b111011101110;
20'b01000100000011110100: color_data = 12'b111011101110;
20'b01000100000011110101: color_data = 12'b111011101110;
20'b01000100000011110110: color_data = 12'b111011101110;
20'b01000100000101001111: color_data = 12'b111011101110;
20'b01000100000101010000: color_data = 12'b111011101110;
20'b01000100000101010001: color_data = 12'b111011101110;
20'b01000100000101010010: color_data = 12'b111011101110;
20'b01000100000101010011: color_data = 12'b111011101110;
20'b01000100000101010100: color_data = 12'b111011101110;
20'b01000100000101010101: color_data = 12'b111011101110;
20'b01000100000101010110: color_data = 12'b111011101110;
20'b01000100000101010111: color_data = 12'b111011101110;
20'b01000100000101011000: color_data = 12'b111011101110;
20'b01000100000110011100: color_data = 12'b111011101110;
20'b01000100000110011101: color_data = 12'b111011101110;
20'b01000100000110011110: color_data = 12'b111011101110;
20'b01000100000110011111: color_data = 12'b111011101110;
20'b01000100000110100000: color_data = 12'b111011101110;
20'b01000100000110100001: color_data = 12'b111011101110;
20'b01000100000110100010: color_data = 12'b111011101110;
20'b01000100000110100011: color_data = 12'b111011101110;
20'b01000100000110100100: color_data = 12'b111011101110;
20'b01000100000110100101: color_data = 12'b111011101110;
20'b01000100000110100111: color_data = 12'b111011101110;
20'b01000100000110101000: color_data = 12'b111011101110;
20'b01000100000110101001: color_data = 12'b111011101110;
20'b01000100000110101010: color_data = 12'b111011101110;
20'b01000100000110101011: color_data = 12'b111011101110;
20'b01000100000110101100: color_data = 12'b111011101110;
20'b01000100000110101101: color_data = 12'b111011101110;
20'b01000100000110101110: color_data = 12'b111011101110;
20'b01000100000110101111: color_data = 12'b111011101110;
20'b01000100000110110000: color_data = 12'b111011101110;
20'b01000100010010010110: color_data = 12'b111011101110;
20'b01000100010010010111: color_data = 12'b111011101110;
20'b01000100010010011000: color_data = 12'b111011101110;
20'b01000100010010011001: color_data = 12'b111011101110;
20'b01000100010010011010: color_data = 12'b111011101110;
20'b01000100010010011011: color_data = 12'b111011101110;
20'b01000100010010011100: color_data = 12'b111011101110;
20'b01000100010010011101: color_data = 12'b111011101110;
20'b01000100010010011110: color_data = 12'b111011101110;
20'b01000100010010011111: color_data = 12'b111011101110;
20'b01000100010011001101: color_data = 12'b111011101110;
20'b01000100010011001110: color_data = 12'b111011101110;
20'b01000100010011001111: color_data = 12'b111011101110;
20'b01000100010011010000: color_data = 12'b111011101110;
20'b01000100010011010001: color_data = 12'b111011101110;
20'b01000100010011010010: color_data = 12'b111011101110;
20'b01000100010011010011: color_data = 12'b111011101110;
20'b01000100010011010100: color_data = 12'b111011101110;
20'b01000100010011010101: color_data = 12'b111011101110;
20'b01000100010011010110: color_data = 12'b111011101110;
20'b01000100010011011000: color_data = 12'b111011101110;
20'b01000100010011011001: color_data = 12'b111011101110;
20'b01000100010011011010: color_data = 12'b111011101110;
20'b01000100010011011011: color_data = 12'b111011101110;
20'b01000100010011011100: color_data = 12'b111011101110;
20'b01000100010011011101: color_data = 12'b111011101110;
20'b01000100010011011110: color_data = 12'b111011101110;
20'b01000100010011011111: color_data = 12'b111011101110;
20'b01000100010011100000: color_data = 12'b111011101110;
20'b01000100010011100001: color_data = 12'b111011101110;
20'b01000100010011101101: color_data = 12'b111011101110;
20'b01000100010011101110: color_data = 12'b111011101110;
20'b01000100010011101111: color_data = 12'b111011101110;
20'b01000100010011110000: color_data = 12'b111011101110;
20'b01000100010011110001: color_data = 12'b111011101110;
20'b01000100010011110010: color_data = 12'b111011101110;
20'b01000100010011110011: color_data = 12'b111011101110;
20'b01000100010011110100: color_data = 12'b111011101110;
20'b01000100010011110101: color_data = 12'b111011101110;
20'b01000100010011110110: color_data = 12'b111011101110;
20'b01000100010101001111: color_data = 12'b111011101110;
20'b01000100010101010000: color_data = 12'b111011101110;
20'b01000100010101010001: color_data = 12'b111011101110;
20'b01000100010101010010: color_data = 12'b111011101110;
20'b01000100010101010011: color_data = 12'b111011101110;
20'b01000100010101010100: color_data = 12'b111011101110;
20'b01000100010101010101: color_data = 12'b111011101110;
20'b01000100010101010110: color_data = 12'b111011101110;
20'b01000100010101010111: color_data = 12'b111011101110;
20'b01000100010101011000: color_data = 12'b111011101110;
20'b01000100010110011100: color_data = 12'b111011101110;
20'b01000100010110011101: color_data = 12'b111011101110;
20'b01000100010110011110: color_data = 12'b111011101110;
20'b01000100010110011111: color_data = 12'b111011101110;
20'b01000100010110100000: color_data = 12'b111011101110;
20'b01000100010110100001: color_data = 12'b111011101110;
20'b01000100010110100010: color_data = 12'b111011101110;
20'b01000100010110100011: color_data = 12'b111011101110;
20'b01000100010110100100: color_data = 12'b111011101110;
20'b01000100010110100101: color_data = 12'b111011101110;
20'b01000100010110100111: color_data = 12'b111011101110;
20'b01000100010110101000: color_data = 12'b111011101110;
20'b01000100010110101001: color_data = 12'b111011101110;
20'b01000100010110101010: color_data = 12'b111011101110;
20'b01000100010110101011: color_data = 12'b111011101110;
20'b01000100010110101100: color_data = 12'b111011101110;
20'b01000100010110101101: color_data = 12'b111011101110;
20'b01000100010110101110: color_data = 12'b111011101110;
20'b01000100010110101111: color_data = 12'b111011101110;
20'b01000100010110110000: color_data = 12'b111011101110;
20'b01000100100010010110: color_data = 12'b111011101110;
20'b01000100100010010111: color_data = 12'b111011101110;
20'b01000100100010011000: color_data = 12'b111011101110;
20'b01000100100010011001: color_data = 12'b111011101110;
20'b01000100100010011010: color_data = 12'b111011101110;
20'b01000100100010011011: color_data = 12'b111011101110;
20'b01000100100010011100: color_data = 12'b111011101110;
20'b01000100100010011101: color_data = 12'b111011101110;
20'b01000100100010011110: color_data = 12'b111011101110;
20'b01000100100010011111: color_data = 12'b111011101110;
20'b01000100100011001101: color_data = 12'b111011101110;
20'b01000100100011001110: color_data = 12'b111011101110;
20'b01000100100011001111: color_data = 12'b111011101110;
20'b01000100100011010000: color_data = 12'b111011101110;
20'b01000100100011010001: color_data = 12'b111011101110;
20'b01000100100011010010: color_data = 12'b111011101110;
20'b01000100100011010011: color_data = 12'b111011101110;
20'b01000100100011010100: color_data = 12'b111011101110;
20'b01000100100011010101: color_data = 12'b111011101110;
20'b01000100100011010110: color_data = 12'b111011101110;
20'b01000100100011011000: color_data = 12'b111011101110;
20'b01000100100011011001: color_data = 12'b111011101110;
20'b01000100100011011010: color_data = 12'b111011101110;
20'b01000100100011011011: color_data = 12'b111011101110;
20'b01000100100011011100: color_data = 12'b111011101110;
20'b01000100100011011101: color_data = 12'b111011101110;
20'b01000100100011011110: color_data = 12'b111011101110;
20'b01000100100011011111: color_data = 12'b111011101110;
20'b01000100100011100000: color_data = 12'b111011101110;
20'b01000100100011100001: color_data = 12'b111011101110;
20'b01000100100011101101: color_data = 12'b111011101110;
20'b01000100100011101110: color_data = 12'b111011101110;
20'b01000100100011101111: color_data = 12'b111011101110;
20'b01000100100011110000: color_data = 12'b111011101110;
20'b01000100100011110001: color_data = 12'b111011101110;
20'b01000100100011110010: color_data = 12'b111011101110;
20'b01000100100011110011: color_data = 12'b111011101110;
20'b01000100100011110100: color_data = 12'b111011101110;
20'b01000100100011110101: color_data = 12'b111011101110;
20'b01000100100011110110: color_data = 12'b111011101110;
20'b01000100100101001111: color_data = 12'b111011101110;
20'b01000100100101010000: color_data = 12'b111011101110;
20'b01000100100101010001: color_data = 12'b111011101110;
20'b01000100100101010010: color_data = 12'b111011101110;
20'b01000100100101010011: color_data = 12'b111011101110;
20'b01000100100101010100: color_data = 12'b111011101110;
20'b01000100100101010101: color_data = 12'b111011101110;
20'b01000100100101010110: color_data = 12'b111011101110;
20'b01000100100101010111: color_data = 12'b111011101110;
20'b01000100100101011000: color_data = 12'b111011101110;
20'b01000100100110011100: color_data = 12'b111011101110;
20'b01000100100110011101: color_data = 12'b111011101110;
20'b01000100100110011110: color_data = 12'b111011101110;
20'b01000100100110011111: color_data = 12'b111011101110;
20'b01000100100110100000: color_data = 12'b111011101110;
20'b01000100100110100001: color_data = 12'b111011101110;
20'b01000100100110100010: color_data = 12'b111011101110;
20'b01000100100110100011: color_data = 12'b111011101110;
20'b01000100100110100100: color_data = 12'b111011101110;
20'b01000100100110100101: color_data = 12'b111011101110;
20'b01000100100110100111: color_data = 12'b111011101110;
20'b01000100100110101000: color_data = 12'b111011101110;
20'b01000100100110101001: color_data = 12'b111011101110;
20'b01000100100110101010: color_data = 12'b111011101110;
20'b01000100100110101011: color_data = 12'b111011101110;
20'b01000100100110101100: color_data = 12'b111011101110;
20'b01000100100110101101: color_data = 12'b111011101110;
20'b01000100100110101110: color_data = 12'b111011101110;
20'b01000100100110101111: color_data = 12'b111011101110;
20'b01000100100110110000: color_data = 12'b111011101110;
20'b01000100110010010110: color_data = 12'b111011101110;
20'b01000100110010010111: color_data = 12'b111011101110;
20'b01000100110010011000: color_data = 12'b111011101110;
20'b01000100110010011001: color_data = 12'b111011101110;
20'b01000100110010011010: color_data = 12'b111011101110;
20'b01000100110010011011: color_data = 12'b111011101110;
20'b01000100110010011100: color_data = 12'b111011101110;
20'b01000100110010011101: color_data = 12'b111011101110;
20'b01000100110010011110: color_data = 12'b111011101110;
20'b01000100110010011111: color_data = 12'b111011101110;
20'b01000100110011001101: color_data = 12'b111011101110;
20'b01000100110011001110: color_data = 12'b111011101110;
20'b01000100110011001111: color_data = 12'b111011101110;
20'b01000100110011010000: color_data = 12'b111011101110;
20'b01000100110011010001: color_data = 12'b111011101110;
20'b01000100110011010010: color_data = 12'b111011101110;
20'b01000100110011010011: color_data = 12'b111011101110;
20'b01000100110011010100: color_data = 12'b111011101110;
20'b01000100110011010101: color_data = 12'b111011101110;
20'b01000100110011010110: color_data = 12'b111011101110;
20'b01000100110011011000: color_data = 12'b111011101110;
20'b01000100110011011001: color_data = 12'b111011101110;
20'b01000100110011011010: color_data = 12'b111011101110;
20'b01000100110011011011: color_data = 12'b111011101110;
20'b01000100110011011100: color_data = 12'b111011101110;
20'b01000100110011011101: color_data = 12'b111011101110;
20'b01000100110011011110: color_data = 12'b111011101110;
20'b01000100110011011111: color_data = 12'b111011101110;
20'b01000100110011100000: color_data = 12'b111011101110;
20'b01000100110011100001: color_data = 12'b111011101110;
20'b01000100110011101101: color_data = 12'b111011101110;
20'b01000100110011101110: color_data = 12'b111011101110;
20'b01000100110011101111: color_data = 12'b111011101110;
20'b01000100110011110000: color_data = 12'b111011101110;
20'b01000100110011110001: color_data = 12'b111011101110;
20'b01000100110011110010: color_data = 12'b111011101110;
20'b01000100110011110011: color_data = 12'b111011101110;
20'b01000100110011110100: color_data = 12'b111011101110;
20'b01000100110011110101: color_data = 12'b111011101110;
20'b01000100110011110110: color_data = 12'b111011101110;
20'b01000100110101001111: color_data = 12'b111011101110;
20'b01000100110101010000: color_data = 12'b111011101110;
20'b01000100110101010001: color_data = 12'b111011101110;
20'b01000100110101010010: color_data = 12'b111011101110;
20'b01000100110101010011: color_data = 12'b111011101110;
20'b01000100110101010100: color_data = 12'b111011101110;
20'b01000100110101010101: color_data = 12'b111011101110;
20'b01000100110101010110: color_data = 12'b111011101110;
20'b01000100110101010111: color_data = 12'b111011101110;
20'b01000100110101011000: color_data = 12'b111011101110;
20'b01000100110110011100: color_data = 12'b111011101110;
20'b01000100110110011101: color_data = 12'b111011101110;
20'b01000100110110011110: color_data = 12'b111011101110;
20'b01000100110110011111: color_data = 12'b111011101110;
20'b01000100110110100000: color_data = 12'b111011101110;
20'b01000100110110100001: color_data = 12'b111011101110;
20'b01000100110110100010: color_data = 12'b111011101110;
20'b01000100110110100011: color_data = 12'b111011101110;
20'b01000100110110100100: color_data = 12'b111011101110;
20'b01000100110110100101: color_data = 12'b111011101110;
20'b01000100110110100111: color_data = 12'b111011101110;
20'b01000100110110101000: color_data = 12'b111011101110;
20'b01000100110110101001: color_data = 12'b111011101110;
20'b01000100110110101010: color_data = 12'b111011101110;
20'b01000100110110101011: color_data = 12'b111011101110;
20'b01000100110110101100: color_data = 12'b111011101110;
20'b01000100110110101101: color_data = 12'b111011101110;
20'b01000100110110101110: color_data = 12'b111011101110;
20'b01000100110110101111: color_data = 12'b111011101110;
20'b01000100110110110000: color_data = 12'b111011101110;
20'b01000101000010010110: color_data = 12'b111011101110;
20'b01000101000010010111: color_data = 12'b111011101110;
20'b01000101000010011000: color_data = 12'b111011101110;
20'b01000101000010011001: color_data = 12'b111011101110;
20'b01000101000010011010: color_data = 12'b111011101110;
20'b01000101000010011011: color_data = 12'b111011101110;
20'b01000101000010011100: color_data = 12'b111011101110;
20'b01000101000010011101: color_data = 12'b111011101110;
20'b01000101000010011110: color_data = 12'b111011101110;
20'b01000101000010011111: color_data = 12'b111011101110;
20'b01000101000011001101: color_data = 12'b111011101110;
20'b01000101000011001110: color_data = 12'b111011101110;
20'b01000101000011001111: color_data = 12'b111011101110;
20'b01000101000011010000: color_data = 12'b111011101110;
20'b01000101000011010001: color_data = 12'b111011101110;
20'b01000101000011010010: color_data = 12'b111011101110;
20'b01000101000011010011: color_data = 12'b111011101110;
20'b01000101000011010100: color_data = 12'b111011101110;
20'b01000101000011010101: color_data = 12'b111011101110;
20'b01000101000011010110: color_data = 12'b111011101110;
20'b01000101000011011000: color_data = 12'b111011101110;
20'b01000101000011011001: color_data = 12'b111011101110;
20'b01000101000011011010: color_data = 12'b111011101110;
20'b01000101000011011011: color_data = 12'b111011101110;
20'b01000101000011011100: color_data = 12'b111011101110;
20'b01000101000011011101: color_data = 12'b111011101110;
20'b01000101000011011110: color_data = 12'b111011101110;
20'b01000101000011011111: color_data = 12'b111011101110;
20'b01000101000011100000: color_data = 12'b111011101110;
20'b01000101000011100001: color_data = 12'b111011101110;
20'b01000101000011101101: color_data = 12'b111011101110;
20'b01000101000011101110: color_data = 12'b111011101110;
20'b01000101000011101111: color_data = 12'b111011101110;
20'b01000101000011110000: color_data = 12'b111011101110;
20'b01000101000011110001: color_data = 12'b111011101110;
20'b01000101000011110010: color_data = 12'b111011101110;
20'b01000101000011110011: color_data = 12'b111011101110;
20'b01000101000011110100: color_data = 12'b111011101110;
20'b01000101000011110101: color_data = 12'b111011101110;
20'b01000101000011110110: color_data = 12'b111011101110;
20'b01000101000101001111: color_data = 12'b111011101110;
20'b01000101000101010000: color_data = 12'b111011101110;
20'b01000101000101010001: color_data = 12'b111011101110;
20'b01000101000101010010: color_data = 12'b111011101110;
20'b01000101000101010011: color_data = 12'b111011101110;
20'b01000101000101010100: color_data = 12'b111011101110;
20'b01000101000101010101: color_data = 12'b111011101110;
20'b01000101000101010110: color_data = 12'b111011101110;
20'b01000101000101010111: color_data = 12'b111011101110;
20'b01000101000101011000: color_data = 12'b111011101110;
20'b01000101000110011100: color_data = 12'b111011101110;
20'b01000101000110011101: color_data = 12'b111011101110;
20'b01000101000110011110: color_data = 12'b111011101110;
20'b01000101000110011111: color_data = 12'b111011101110;
20'b01000101000110100000: color_data = 12'b111011101110;
20'b01000101000110100001: color_data = 12'b111011101110;
20'b01000101000110100010: color_data = 12'b111011101110;
20'b01000101000110100011: color_data = 12'b111011101110;
20'b01000101000110100100: color_data = 12'b111011101110;
20'b01000101000110100101: color_data = 12'b111011101110;
20'b01000101000110100111: color_data = 12'b111011101110;
20'b01000101000110101000: color_data = 12'b111011101110;
20'b01000101000110101001: color_data = 12'b111011101110;
20'b01000101000110101010: color_data = 12'b111011101110;
20'b01000101000110101011: color_data = 12'b111011101110;
20'b01000101000110101100: color_data = 12'b111011101110;
20'b01000101000110101101: color_data = 12'b111011101110;
20'b01000101000110101110: color_data = 12'b111011101110;
20'b01000101000110101111: color_data = 12'b111011101110;
20'b01000101000110110000: color_data = 12'b111011101110;
20'b01000101100010010110: color_data = 12'b111011101110;
20'b01000101100010010111: color_data = 12'b111011101110;
20'b01000101100010011000: color_data = 12'b111011101110;
20'b01000101100010011001: color_data = 12'b111011101110;
20'b01000101100010011010: color_data = 12'b111011101110;
20'b01000101100010011011: color_data = 12'b111011101110;
20'b01000101100010011100: color_data = 12'b111011101110;
20'b01000101100010011101: color_data = 12'b111011101110;
20'b01000101100010011110: color_data = 12'b111011101110;
20'b01000101100010011111: color_data = 12'b111011101110;
20'b01000101100010100001: color_data = 12'b111011101110;
20'b01000101100010100010: color_data = 12'b111011101110;
20'b01000101100010100011: color_data = 12'b111011101110;
20'b01000101100010100100: color_data = 12'b111011101110;
20'b01000101100010100101: color_data = 12'b111011101110;
20'b01000101100010100110: color_data = 12'b111011101110;
20'b01000101100010100111: color_data = 12'b111011101110;
20'b01000101100010101000: color_data = 12'b111011101110;
20'b01000101100010101001: color_data = 12'b111011101110;
20'b01000101100010101010: color_data = 12'b111011101110;
20'b01000101100011001101: color_data = 12'b111011101110;
20'b01000101100011001110: color_data = 12'b111011101110;
20'b01000101100011001111: color_data = 12'b111011101110;
20'b01000101100011010000: color_data = 12'b111011101110;
20'b01000101100011010001: color_data = 12'b111011101110;
20'b01000101100011010010: color_data = 12'b111011101110;
20'b01000101100011010011: color_data = 12'b111011101110;
20'b01000101100011010100: color_data = 12'b111011101110;
20'b01000101100011010101: color_data = 12'b111011101110;
20'b01000101100011010110: color_data = 12'b111011101110;
20'b01000101100011011000: color_data = 12'b111011101110;
20'b01000101100011011001: color_data = 12'b111011101110;
20'b01000101100011011010: color_data = 12'b111011101110;
20'b01000101100011011011: color_data = 12'b111011101110;
20'b01000101100011011100: color_data = 12'b111011101110;
20'b01000101100011011101: color_data = 12'b111011101110;
20'b01000101100011011110: color_data = 12'b111011101110;
20'b01000101100011011111: color_data = 12'b111011101110;
20'b01000101100011100000: color_data = 12'b111011101110;
20'b01000101100011100001: color_data = 12'b111011101110;
20'b01000101100011101101: color_data = 12'b111011101110;
20'b01000101100011101110: color_data = 12'b111011101110;
20'b01000101100011101111: color_data = 12'b111011101110;
20'b01000101100011110000: color_data = 12'b111011101110;
20'b01000101100011110001: color_data = 12'b111011101110;
20'b01000101100011110010: color_data = 12'b111011101110;
20'b01000101100011110011: color_data = 12'b111011101110;
20'b01000101100011110100: color_data = 12'b111011101110;
20'b01000101100011110101: color_data = 12'b111011101110;
20'b01000101100011110110: color_data = 12'b111011101110;
20'b01000101100011111000: color_data = 12'b111011101110;
20'b01000101100011111001: color_data = 12'b111011101110;
20'b01000101100011111010: color_data = 12'b111011101110;
20'b01000101100011111011: color_data = 12'b111011101110;
20'b01000101100011111100: color_data = 12'b111011101110;
20'b01000101100011111101: color_data = 12'b111011101110;
20'b01000101100011111110: color_data = 12'b111011101110;
20'b01000101100011111111: color_data = 12'b111011101110;
20'b01000101100100000000: color_data = 12'b111011101110;
20'b01000101100100000001: color_data = 12'b111011101110;
20'b01000101100100100100: color_data = 12'b111011101110;
20'b01000101100100100101: color_data = 12'b111011101110;
20'b01000101100100100110: color_data = 12'b111011101110;
20'b01000101100100100111: color_data = 12'b111011101110;
20'b01000101100100101000: color_data = 12'b111011101110;
20'b01000101100100101001: color_data = 12'b111011101110;
20'b01000101100100101010: color_data = 12'b111011101110;
20'b01000101100100101011: color_data = 12'b111011101110;
20'b01000101100100101100: color_data = 12'b111011101110;
20'b01000101100100101101: color_data = 12'b111011101110;
20'b01000101100100101111: color_data = 12'b111011101110;
20'b01000101100100110000: color_data = 12'b111011101110;
20'b01000101100100110001: color_data = 12'b111011101110;
20'b01000101100100110010: color_data = 12'b111011101110;
20'b01000101100100110011: color_data = 12'b111011101110;
20'b01000101100100110100: color_data = 12'b111011101110;
20'b01000101100100110101: color_data = 12'b111011101110;
20'b01000101100100110110: color_data = 12'b111011101110;
20'b01000101100100110111: color_data = 12'b111011101110;
20'b01000101100100111000: color_data = 12'b111011101110;
20'b01000101100101000100: color_data = 12'b111011101110;
20'b01000101100101000101: color_data = 12'b111011101110;
20'b01000101100101000110: color_data = 12'b111011101110;
20'b01000101100101000111: color_data = 12'b111011101110;
20'b01000101100101001000: color_data = 12'b111011101110;
20'b01000101100101001001: color_data = 12'b111011101110;
20'b01000101100101001010: color_data = 12'b111011101110;
20'b01000101100101001011: color_data = 12'b111011101110;
20'b01000101100101001100: color_data = 12'b111011101110;
20'b01000101100101001101: color_data = 12'b111011101110;
20'b01000101100101001111: color_data = 12'b111011101110;
20'b01000101100101010000: color_data = 12'b111011101110;
20'b01000101100101010001: color_data = 12'b111011101110;
20'b01000101100101010010: color_data = 12'b111011101110;
20'b01000101100101010011: color_data = 12'b111011101110;
20'b01000101100101010100: color_data = 12'b111011101110;
20'b01000101100101010101: color_data = 12'b111011101110;
20'b01000101100101010110: color_data = 12'b111011101110;
20'b01000101100101010111: color_data = 12'b111011101110;
20'b01000101100101011000: color_data = 12'b111011101110;
20'b01000101100110011100: color_data = 12'b111011101110;
20'b01000101100110011101: color_data = 12'b111011101110;
20'b01000101100110011110: color_data = 12'b111011101110;
20'b01000101100110011111: color_data = 12'b111011101110;
20'b01000101100110100000: color_data = 12'b111011101110;
20'b01000101100110100001: color_data = 12'b111011101110;
20'b01000101100110100010: color_data = 12'b111011101110;
20'b01000101100110100011: color_data = 12'b111011101110;
20'b01000101100110100100: color_data = 12'b111011101110;
20'b01000101100110100101: color_data = 12'b111011101110;
20'b01000101100110100111: color_data = 12'b111011101110;
20'b01000101100110101000: color_data = 12'b111011101110;
20'b01000101100110101001: color_data = 12'b111011101110;
20'b01000101100110101010: color_data = 12'b111011101110;
20'b01000101100110101011: color_data = 12'b111011101110;
20'b01000101100110101100: color_data = 12'b111011101110;
20'b01000101100110101101: color_data = 12'b111011101110;
20'b01000101100110101110: color_data = 12'b111011101110;
20'b01000101100110101111: color_data = 12'b111011101110;
20'b01000101100110110000: color_data = 12'b111011101110;
20'b01000101100111010011: color_data = 12'b111011101110;
20'b01000101100111010100: color_data = 12'b111011101110;
20'b01000101100111010101: color_data = 12'b111011101110;
20'b01000101100111010110: color_data = 12'b111011101110;
20'b01000101100111010111: color_data = 12'b111011101110;
20'b01000101100111011000: color_data = 12'b111011101110;
20'b01000101100111011001: color_data = 12'b111011101110;
20'b01000101100111011010: color_data = 12'b111011101110;
20'b01000101100111011011: color_data = 12'b111011101110;
20'b01000101100111011100: color_data = 12'b111011101110;
20'b01000101100111011110: color_data = 12'b111011101110;
20'b01000101100111011111: color_data = 12'b111011101110;
20'b01000101100111100000: color_data = 12'b111011101110;
20'b01000101100111100001: color_data = 12'b111011101110;
20'b01000101100111100010: color_data = 12'b111011101110;
20'b01000101100111100011: color_data = 12'b111011101110;
20'b01000101100111100100: color_data = 12'b111011101110;
20'b01000101100111100101: color_data = 12'b111011101110;
20'b01000101100111100110: color_data = 12'b111011101110;
20'b01000101100111100111: color_data = 12'b111011101110;
20'b01000101110010010110: color_data = 12'b111011101110;
20'b01000101110010010111: color_data = 12'b111011101110;
20'b01000101110010011000: color_data = 12'b111011101110;
20'b01000101110010011001: color_data = 12'b111011101110;
20'b01000101110010011010: color_data = 12'b111011101110;
20'b01000101110010011011: color_data = 12'b111011101110;
20'b01000101110010011100: color_data = 12'b111011101110;
20'b01000101110010011101: color_data = 12'b111011101110;
20'b01000101110010011110: color_data = 12'b111011101110;
20'b01000101110010011111: color_data = 12'b111011101110;
20'b01000101110010100001: color_data = 12'b111011101110;
20'b01000101110010100010: color_data = 12'b111011101110;
20'b01000101110010100011: color_data = 12'b111011101110;
20'b01000101110010100100: color_data = 12'b111011101110;
20'b01000101110010100101: color_data = 12'b111011101110;
20'b01000101110010100110: color_data = 12'b111011101110;
20'b01000101110010100111: color_data = 12'b111011101110;
20'b01000101110010101000: color_data = 12'b111011101110;
20'b01000101110010101001: color_data = 12'b111011101110;
20'b01000101110010101010: color_data = 12'b111011101110;
20'b01000101110011001101: color_data = 12'b111011101110;
20'b01000101110011001110: color_data = 12'b111011101110;
20'b01000101110011001111: color_data = 12'b111011101110;
20'b01000101110011010000: color_data = 12'b111011101110;
20'b01000101110011010001: color_data = 12'b111011101110;
20'b01000101110011010010: color_data = 12'b111011101110;
20'b01000101110011010011: color_data = 12'b111011101110;
20'b01000101110011010100: color_data = 12'b111011101110;
20'b01000101110011010101: color_data = 12'b111011101110;
20'b01000101110011010110: color_data = 12'b111011101110;
20'b01000101110011011000: color_data = 12'b111011101110;
20'b01000101110011011001: color_data = 12'b111011101110;
20'b01000101110011011010: color_data = 12'b111011101110;
20'b01000101110011011011: color_data = 12'b111011101110;
20'b01000101110011011100: color_data = 12'b111011101110;
20'b01000101110011011101: color_data = 12'b111011101110;
20'b01000101110011011110: color_data = 12'b111011101110;
20'b01000101110011011111: color_data = 12'b111011101110;
20'b01000101110011100000: color_data = 12'b111011101110;
20'b01000101110011100001: color_data = 12'b111011101110;
20'b01000101110011101101: color_data = 12'b111011101110;
20'b01000101110011101110: color_data = 12'b111011101110;
20'b01000101110011101111: color_data = 12'b111011101110;
20'b01000101110011110000: color_data = 12'b111011101110;
20'b01000101110011110001: color_data = 12'b111011101110;
20'b01000101110011110010: color_data = 12'b111011101110;
20'b01000101110011110011: color_data = 12'b111011101110;
20'b01000101110011110100: color_data = 12'b111011101110;
20'b01000101110011110101: color_data = 12'b111011101110;
20'b01000101110011110110: color_data = 12'b111011101110;
20'b01000101110011111000: color_data = 12'b111011101110;
20'b01000101110011111001: color_data = 12'b111011101110;
20'b01000101110011111010: color_data = 12'b111011101110;
20'b01000101110011111011: color_data = 12'b111011101110;
20'b01000101110011111100: color_data = 12'b111011101110;
20'b01000101110011111101: color_data = 12'b111011101110;
20'b01000101110011111110: color_data = 12'b111011101110;
20'b01000101110011111111: color_data = 12'b111011101110;
20'b01000101110100000000: color_data = 12'b111011101110;
20'b01000101110100000001: color_data = 12'b111011101110;
20'b01000101110100100100: color_data = 12'b111011101110;
20'b01000101110100100101: color_data = 12'b111011101110;
20'b01000101110100100110: color_data = 12'b111011101110;
20'b01000101110100100111: color_data = 12'b111011101110;
20'b01000101110100101000: color_data = 12'b111011101110;
20'b01000101110100101001: color_data = 12'b111011101110;
20'b01000101110100101010: color_data = 12'b111011101110;
20'b01000101110100101011: color_data = 12'b111011101110;
20'b01000101110100101100: color_data = 12'b111011101110;
20'b01000101110100101101: color_data = 12'b111011101110;
20'b01000101110100101111: color_data = 12'b111011101110;
20'b01000101110100110000: color_data = 12'b111011101110;
20'b01000101110100110001: color_data = 12'b111011101110;
20'b01000101110100110010: color_data = 12'b111011101110;
20'b01000101110100110011: color_data = 12'b111011101110;
20'b01000101110100110100: color_data = 12'b111011101110;
20'b01000101110100110101: color_data = 12'b111011101110;
20'b01000101110100110110: color_data = 12'b111011101110;
20'b01000101110100110111: color_data = 12'b111011101110;
20'b01000101110100111000: color_data = 12'b111011101110;
20'b01000101110101000100: color_data = 12'b111011101110;
20'b01000101110101000101: color_data = 12'b111011101110;
20'b01000101110101000110: color_data = 12'b111011101110;
20'b01000101110101000111: color_data = 12'b111011101110;
20'b01000101110101001000: color_data = 12'b111011101110;
20'b01000101110101001001: color_data = 12'b111011101110;
20'b01000101110101001010: color_data = 12'b111011101110;
20'b01000101110101001011: color_data = 12'b111011101110;
20'b01000101110101001100: color_data = 12'b111011101110;
20'b01000101110101001101: color_data = 12'b111011101110;
20'b01000101110101001111: color_data = 12'b111011101110;
20'b01000101110101010000: color_data = 12'b111011101110;
20'b01000101110101010001: color_data = 12'b111011101110;
20'b01000101110101010010: color_data = 12'b111011101110;
20'b01000101110101010011: color_data = 12'b111011101110;
20'b01000101110101010100: color_data = 12'b111011101110;
20'b01000101110101010101: color_data = 12'b111011101110;
20'b01000101110101010110: color_data = 12'b111011101110;
20'b01000101110101010111: color_data = 12'b111011101110;
20'b01000101110101011000: color_data = 12'b111011101110;
20'b01000101110110011100: color_data = 12'b111011101110;
20'b01000101110110011101: color_data = 12'b111011101110;
20'b01000101110110011110: color_data = 12'b111011101110;
20'b01000101110110011111: color_data = 12'b111011101110;
20'b01000101110110100000: color_data = 12'b111011101110;
20'b01000101110110100001: color_data = 12'b111011101110;
20'b01000101110110100010: color_data = 12'b111011101110;
20'b01000101110110100011: color_data = 12'b111011101110;
20'b01000101110110100100: color_data = 12'b111011101110;
20'b01000101110110100101: color_data = 12'b111011101110;
20'b01000101110110100111: color_data = 12'b111011101110;
20'b01000101110110101000: color_data = 12'b111011101110;
20'b01000101110110101001: color_data = 12'b111011101110;
20'b01000101110110101010: color_data = 12'b111011101110;
20'b01000101110110101011: color_data = 12'b111011101110;
20'b01000101110110101100: color_data = 12'b111011101110;
20'b01000101110110101101: color_data = 12'b111011101110;
20'b01000101110110101110: color_data = 12'b111011101110;
20'b01000101110110101111: color_data = 12'b111011101110;
20'b01000101110110110000: color_data = 12'b111011101110;
20'b01000101110111010011: color_data = 12'b111011101110;
20'b01000101110111010100: color_data = 12'b111011101110;
20'b01000101110111010101: color_data = 12'b111011101110;
20'b01000101110111010110: color_data = 12'b111011101110;
20'b01000101110111010111: color_data = 12'b111011101110;
20'b01000101110111011000: color_data = 12'b111011101110;
20'b01000101110111011001: color_data = 12'b111011101110;
20'b01000101110111011010: color_data = 12'b111011101110;
20'b01000101110111011011: color_data = 12'b111011101110;
20'b01000101110111011100: color_data = 12'b111011101110;
20'b01000101110111011110: color_data = 12'b111011101110;
20'b01000101110111011111: color_data = 12'b111011101110;
20'b01000101110111100000: color_data = 12'b111011101110;
20'b01000101110111100001: color_data = 12'b111011101110;
20'b01000101110111100010: color_data = 12'b111011101110;
20'b01000101110111100011: color_data = 12'b111011101110;
20'b01000101110111100100: color_data = 12'b111011101110;
20'b01000101110111100101: color_data = 12'b111011101110;
20'b01000101110111100110: color_data = 12'b111011101110;
20'b01000101110111100111: color_data = 12'b111011101110;
20'b01000110000010010110: color_data = 12'b111011101110;
20'b01000110000010010111: color_data = 12'b111011101110;
20'b01000110000010011000: color_data = 12'b111011101110;
20'b01000110000010011001: color_data = 12'b111011101110;
20'b01000110000010011010: color_data = 12'b111011101110;
20'b01000110000010011011: color_data = 12'b111011101110;
20'b01000110000010011100: color_data = 12'b111011101110;
20'b01000110000010011101: color_data = 12'b111011101110;
20'b01000110000010011110: color_data = 12'b111011101110;
20'b01000110000010011111: color_data = 12'b111011101110;
20'b01000110000010100001: color_data = 12'b111011101110;
20'b01000110000010100010: color_data = 12'b111011101110;
20'b01000110000010100011: color_data = 12'b111011101110;
20'b01000110000010100100: color_data = 12'b111011101110;
20'b01000110000010100101: color_data = 12'b111011101110;
20'b01000110000010100110: color_data = 12'b111011101110;
20'b01000110000010100111: color_data = 12'b111011101110;
20'b01000110000010101000: color_data = 12'b111011101110;
20'b01000110000010101001: color_data = 12'b111011101110;
20'b01000110000010101010: color_data = 12'b111011101110;
20'b01000110000011001101: color_data = 12'b111011101110;
20'b01000110000011001110: color_data = 12'b111011101110;
20'b01000110000011001111: color_data = 12'b111011101110;
20'b01000110000011010000: color_data = 12'b111011101110;
20'b01000110000011010001: color_data = 12'b111011101110;
20'b01000110000011010010: color_data = 12'b111011101110;
20'b01000110000011010011: color_data = 12'b111011101110;
20'b01000110000011010100: color_data = 12'b111011101110;
20'b01000110000011010101: color_data = 12'b111011101110;
20'b01000110000011010110: color_data = 12'b111011101110;
20'b01000110000011011000: color_data = 12'b111011101110;
20'b01000110000011011001: color_data = 12'b111011101110;
20'b01000110000011011010: color_data = 12'b111011101110;
20'b01000110000011011011: color_data = 12'b111011101110;
20'b01000110000011011100: color_data = 12'b111011101110;
20'b01000110000011011101: color_data = 12'b111011101110;
20'b01000110000011011110: color_data = 12'b111011101110;
20'b01000110000011011111: color_data = 12'b111011101110;
20'b01000110000011100000: color_data = 12'b111011101110;
20'b01000110000011100001: color_data = 12'b111011101110;
20'b01000110000011101101: color_data = 12'b111011101110;
20'b01000110000011101110: color_data = 12'b111011101110;
20'b01000110000011101111: color_data = 12'b111011101110;
20'b01000110000011110000: color_data = 12'b111011101110;
20'b01000110000011110001: color_data = 12'b111011101110;
20'b01000110000011110010: color_data = 12'b111011101110;
20'b01000110000011110011: color_data = 12'b111011101110;
20'b01000110000011110100: color_data = 12'b111011101110;
20'b01000110000011110101: color_data = 12'b111011101110;
20'b01000110000011110110: color_data = 12'b111011101110;
20'b01000110000011111000: color_data = 12'b111011101110;
20'b01000110000011111001: color_data = 12'b111011101110;
20'b01000110000011111010: color_data = 12'b111011101110;
20'b01000110000011111011: color_data = 12'b111011101110;
20'b01000110000011111100: color_data = 12'b111011101110;
20'b01000110000011111101: color_data = 12'b111011101110;
20'b01000110000011111110: color_data = 12'b111011101110;
20'b01000110000011111111: color_data = 12'b111011101110;
20'b01000110000100000000: color_data = 12'b111011101110;
20'b01000110000100000001: color_data = 12'b111011101110;
20'b01000110000100100100: color_data = 12'b111011101110;
20'b01000110000100100101: color_data = 12'b111011101110;
20'b01000110000100100110: color_data = 12'b111011101110;
20'b01000110000100100111: color_data = 12'b111011101110;
20'b01000110000100101000: color_data = 12'b111011101110;
20'b01000110000100101001: color_data = 12'b111011101110;
20'b01000110000100101010: color_data = 12'b111011101110;
20'b01000110000100101011: color_data = 12'b111011101110;
20'b01000110000100101100: color_data = 12'b111011101110;
20'b01000110000100101101: color_data = 12'b111011101110;
20'b01000110000100101111: color_data = 12'b111011101110;
20'b01000110000100110000: color_data = 12'b111011101110;
20'b01000110000100110001: color_data = 12'b111011101110;
20'b01000110000100110010: color_data = 12'b111011101110;
20'b01000110000100110011: color_data = 12'b111011101110;
20'b01000110000100110100: color_data = 12'b111011101110;
20'b01000110000100110101: color_data = 12'b111011101110;
20'b01000110000100110110: color_data = 12'b111011101110;
20'b01000110000100110111: color_data = 12'b111011101110;
20'b01000110000100111000: color_data = 12'b111011101110;
20'b01000110000101000100: color_data = 12'b111011101110;
20'b01000110000101000101: color_data = 12'b111011101110;
20'b01000110000101000110: color_data = 12'b111011101110;
20'b01000110000101000111: color_data = 12'b111011101110;
20'b01000110000101001000: color_data = 12'b111011101110;
20'b01000110000101001001: color_data = 12'b111011101110;
20'b01000110000101001010: color_data = 12'b111011101110;
20'b01000110000101001011: color_data = 12'b111011101110;
20'b01000110000101001100: color_data = 12'b111011101110;
20'b01000110000101001101: color_data = 12'b111011101110;
20'b01000110000101001111: color_data = 12'b111011101110;
20'b01000110000101010000: color_data = 12'b111011101110;
20'b01000110000101010001: color_data = 12'b111011101110;
20'b01000110000101010010: color_data = 12'b111011101110;
20'b01000110000101010011: color_data = 12'b111011101110;
20'b01000110000101010100: color_data = 12'b111011101110;
20'b01000110000101010101: color_data = 12'b111011101110;
20'b01000110000101010110: color_data = 12'b111011101110;
20'b01000110000101010111: color_data = 12'b111011101110;
20'b01000110000101011000: color_data = 12'b111011101110;
20'b01000110000110011100: color_data = 12'b111011101110;
20'b01000110000110011101: color_data = 12'b111011101110;
20'b01000110000110011110: color_data = 12'b111011101110;
20'b01000110000110011111: color_data = 12'b111011101110;
20'b01000110000110100000: color_data = 12'b111011101110;
20'b01000110000110100001: color_data = 12'b111011101110;
20'b01000110000110100010: color_data = 12'b111011101110;
20'b01000110000110100011: color_data = 12'b111011101110;
20'b01000110000110100100: color_data = 12'b111011101110;
20'b01000110000110100101: color_data = 12'b111011101110;
20'b01000110000110100111: color_data = 12'b111011101110;
20'b01000110000110101000: color_data = 12'b111011101110;
20'b01000110000110101001: color_data = 12'b111011101110;
20'b01000110000110101010: color_data = 12'b111011101110;
20'b01000110000110101011: color_data = 12'b111011101110;
20'b01000110000110101100: color_data = 12'b111011101110;
20'b01000110000110101101: color_data = 12'b111011101110;
20'b01000110000110101110: color_data = 12'b111011101110;
20'b01000110000110101111: color_data = 12'b111011101110;
20'b01000110000110110000: color_data = 12'b111011101110;
20'b01000110000111010011: color_data = 12'b111011101110;
20'b01000110000111010100: color_data = 12'b111011101110;
20'b01000110000111010101: color_data = 12'b111011101110;
20'b01000110000111010110: color_data = 12'b111011101110;
20'b01000110000111010111: color_data = 12'b111011101110;
20'b01000110000111011000: color_data = 12'b111011101110;
20'b01000110000111011001: color_data = 12'b111011101110;
20'b01000110000111011010: color_data = 12'b111011101110;
20'b01000110000111011011: color_data = 12'b111011101110;
20'b01000110000111011100: color_data = 12'b111011101110;
20'b01000110000111011110: color_data = 12'b111011101110;
20'b01000110000111011111: color_data = 12'b111011101110;
20'b01000110000111100000: color_data = 12'b111011101110;
20'b01000110000111100001: color_data = 12'b111011101110;
20'b01000110000111100010: color_data = 12'b111011101110;
20'b01000110000111100011: color_data = 12'b111011101110;
20'b01000110000111100100: color_data = 12'b111011101110;
20'b01000110000111100101: color_data = 12'b111011101110;
20'b01000110000111100110: color_data = 12'b111011101110;
20'b01000110000111100111: color_data = 12'b111011101110;
20'b01000110010010010110: color_data = 12'b111011101110;
20'b01000110010010010111: color_data = 12'b111011101110;
20'b01000110010010011000: color_data = 12'b111011101110;
20'b01000110010010011001: color_data = 12'b111011101110;
20'b01000110010010011010: color_data = 12'b111011101110;
20'b01000110010010011011: color_data = 12'b111011101110;
20'b01000110010010011100: color_data = 12'b111011101110;
20'b01000110010010011101: color_data = 12'b111011101110;
20'b01000110010010011110: color_data = 12'b111011101110;
20'b01000110010010011111: color_data = 12'b111011101110;
20'b01000110010010100001: color_data = 12'b111011101110;
20'b01000110010010100010: color_data = 12'b111011101110;
20'b01000110010010100011: color_data = 12'b111011101110;
20'b01000110010010100100: color_data = 12'b111011101110;
20'b01000110010010100101: color_data = 12'b111011101110;
20'b01000110010010100110: color_data = 12'b111011101110;
20'b01000110010010100111: color_data = 12'b111011101110;
20'b01000110010010101000: color_data = 12'b111011101110;
20'b01000110010010101001: color_data = 12'b111011101110;
20'b01000110010010101010: color_data = 12'b111011101110;
20'b01000110010011001101: color_data = 12'b111011101110;
20'b01000110010011001110: color_data = 12'b111011101110;
20'b01000110010011001111: color_data = 12'b111011101110;
20'b01000110010011010000: color_data = 12'b111011101110;
20'b01000110010011010001: color_data = 12'b111011101110;
20'b01000110010011010010: color_data = 12'b111011101110;
20'b01000110010011010011: color_data = 12'b111011101110;
20'b01000110010011010100: color_data = 12'b111011101110;
20'b01000110010011010101: color_data = 12'b111011101110;
20'b01000110010011010110: color_data = 12'b111011101110;
20'b01000110010011011000: color_data = 12'b111011101110;
20'b01000110010011011001: color_data = 12'b111011101110;
20'b01000110010011011010: color_data = 12'b111011101110;
20'b01000110010011011011: color_data = 12'b111011101110;
20'b01000110010011011100: color_data = 12'b111011101110;
20'b01000110010011011101: color_data = 12'b111011101110;
20'b01000110010011011110: color_data = 12'b111011101110;
20'b01000110010011011111: color_data = 12'b111011101110;
20'b01000110010011100000: color_data = 12'b111011101110;
20'b01000110010011100001: color_data = 12'b111011101110;
20'b01000110010011101101: color_data = 12'b111011101110;
20'b01000110010011101110: color_data = 12'b111011101110;
20'b01000110010011101111: color_data = 12'b111011101110;
20'b01000110010011110000: color_data = 12'b111011101110;
20'b01000110010011110001: color_data = 12'b111011101110;
20'b01000110010011110010: color_data = 12'b111011101110;
20'b01000110010011110011: color_data = 12'b111011101110;
20'b01000110010011110100: color_data = 12'b111011101110;
20'b01000110010011110101: color_data = 12'b111011101110;
20'b01000110010011110110: color_data = 12'b111011101110;
20'b01000110010011111000: color_data = 12'b111011101110;
20'b01000110010011111001: color_data = 12'b111011101110;
20'b01000110010011111010: color_data = 12'b111011101110;
20'b01000110010011111011: color_data = 12'b111011101110;
20'b01000110010011111100: color_data = 12'b111011101110;
20'b01000110010011111101: color_data = 12'b111011101110;
20'b01000110010011111110: color_data = 12'b111011101110;
20'b01000110010011111111: color_data = 12'b111011101110;
20'b01000110010100000000: color_data = 12'b111011101110;
20'b01000110010100000001: color_data = 12'b111011101110;
20'b01000110010100100100: color_data = 12'b111011101110;
20'b01000110010100100101: color_data = 12'b111011101110;
20'b01000110010100100110: color_data = 12'b111011101110;
20'b01000110010100100111: color_data = 12'b111011101110;
20'b01000110010100101000: color_data = 12'b111011101110;
20'b01000110010100101001: color_data = 12'b111011101110;
20'b01000110010100101010: color_data = 12'b111011101110;
20'b01000110010100101011: color_data = 12'b111011101110;
20'b01000110010100101100: color_data = 12'b111011101110;
20'b01000110010100101101: color_data = 12'b111011101110;
20'b01000110010100101111: color_data = 12'b111011101110;
20'b01000110010100110000: color_data = 12'b111011101110;
20'b01000110010100110001: color_data = 12'b111011101110;
20'b01000110010100110010: color_data = 12'b111011101110;
20'b01000110010100110011: color_data = 12'b111011101110;
20'b01000110010100110100: color_data = 12'b111011101110;
20'b01000110010100110101: color_data = 12'b111011101110;
20'b01000110010100110110: color_data = 12'b111011101110;
20'b01000110010100110111: color_data = 12'b111011101110;
20'b01000110010100111000: color_data = 12'b111011101110;
20'b01000110010101000100: color_data = 12'b111011101110;
20'b01000110010101000101: color_data = 12'b111011101110;
20'b01000110010101000110: color_data = 12'b111011101110;
20'b01000110010101000111: color_data = 12'b111011101110;
20'b01000110010101001000: color_data = 12'b111011101110;
20'b01000110010101001001: color_data = 12'b111011101110;
20'b01000110010101001010: color_data = 12'b111011101110;
20'b01000110010101001011: color_data = 12'b111011101110;
20'b01000110010101001100: color_data = 12'b111011101110;
20'b01000110010101001101: color_data = 12'b111011101110;
20'b01000110010101001111: color_data = 12'b111011101110;
20'b01000110010101010000: color_data = 12'b111011101110;
20'b01000110010101010001: color_data = 12'b111011101110;
20'b01000110010101010010: color_data = 12'b111011101110;
20'b01000110010101010011: color_data = 12'b111011101110;
20'b01000110010101010100: color_data = 12'b111011101110;
20'b01000110010101010101: color_data = 12'b111011101110;
20'b01000110010101010110: color_data = 12'b111011101110;
20'b01000110010101010111: color_data = 12'b111011101110;
20'b01000110010101011000: color_data = 12'b111011101110;
20'b01000110010110011100: color_data = 12'b111011101110;
20'b01000110010110011101: color_data = 12'b111011101110;
20'b01000110010110011110: color_data = 12'b111011101110;
20'b01000110010110011111: color_data = 12'b111011101110;
20'b01000110010110100000: color_data = 12'b111011101110;
20'b01000110010110100001: color_data = 12'b111011101110;
20'b01000110010110100010: color_data = 12'b111011101110;
20'b01000110010110100011: color_data = 12'b111011101110;
20'b01000110010110100100: color_data = 12'b111011101110;
20'b01000110010110100101: color_data = 12'b111011101110;
20'b01000110010110100111: color_data = 12'b111011101110;
20'b01000110010110101000: color_data = 12'b111011101110;
20'b01000110010110101001: color_data = 12'b111011101110;
20'b01000110010110101010: color_data = 12'b111011101110;
20'b01000110010110101011: color_data = 12'b111011101110;
20'b01000110010110101100: color_data = 12'b111011101110;
20'b01000110010110101101: color_data = 12'b111011101110;
20'b01000110010110101110: color_data = 12'b111011101110;
20'b01000110010110101111: color_data = 12'b111011101110;
20'b01000110010110110000: color_data = 12'b111011101110;
20'b01000110010111010011: color_data = 12'b111011101110;
20'b01000110010111010100: color_data = 12'b111011101110;
20'b01000110010111010101: color_data = 12'b111011101110;
20'b01000110010111010110: color_data = 12'b111011101110;
20'b01000110010111010111: color_data = 12'b111011101110;
20'b01000110010111011000: color_data = 12'b111011101110;
20'b01000110010111011001: color_data = 12'b111011101110;
20'b01000110010111011010: color_data = 12'b111011101110;
20'b01000110010111011011: color_data = 12'b111011101110;
20'b01000110010111011100: color_data = 12'b111011101110;
20'b01000110010111011110: color_data = 12'b111011101110;
20'b01000110010111011111: color_data = 12'b111011101110;
20'b01000110010111100000: color_data = 12'b111011101110;
20'b01000110010111100001: color_data = 12'b111011101110;
20'b01000110010111100010: color_data = 12'b111011101110;
20'b01000110010111100011: color_data = 12'b111011101110;
20'b01000110010111100100: color_data = 12'b111011101110;
20'b01000110010111100101: color_data = 12'b111011101110;
20'b01000110010111100110: color_data = 12'b111011101110;
20'b01000110010111100111: color_data = 12'b111011101110;
20'b01000110100010010110: color_data = 12'b111011101110;
20'b01000110100010010111: color_data = 12'b111011101110;
20'b01000110100010011000: color_data = 12'b111011101110;
20'b01000110100010011001: color_data = 12'b111011101110;
20'b01000110100010011010: color_data = 12'b111011101110;
20'b01000110100010011011: color_data = 12'b111011101110;
20'b01000110100010011100: color_data = 12'b111011101110;
20'b01000110100010011101: color_data = 12'b111011101110;
20'b01000110100010011110: color_data = 12'b111011101110;
20'b01000110100010011111: color_data = 12'b111011101110;
20'b01000110100010100001: color_data = 12'b111011101110;
20'b01000110100010100010: color_data = 12'b111011101110;
20'b01000110100010100011: color_data = 12'b111011101110;
20'b01000110100010100100: color_data = 12'b111011101110;
20'b01000110100010100101: color_data = 12'b111011101110;
20'b01000110100010100110: color_data = 12'b111011101110;
20'b01000110100010100111: color_data = 12'b111011101110;
20'b01000110100010101000: color_data = 12'b111011101110;
20'b01000110100010101001: color_data = 12'b111011101110;
20'b01000110100010101010: color_data = 12'b111011101110;
20'b01000110100011001101: color_data = 12'b111011101110;
20'b01000110100011001110: color_data = 12'b111011101110;
20'b01000110100011001111: color_data = 12'b111011101110;
20'b01000110100011010000: color_data = 12'b111011101110;
20'b01000110100011010001: color_data = 12'b111011101110;
20'b01000110100011010010: color_data = 12'b111011101110;
20'b01000110100011010011: color_data = 12'b111011101110;
20'b01000110100011010100: color_data = 12'b111011101110;
20'b01000110100011010101: color_data = 12'b111011101110;
20'b01000110100011010110: color_data = 12'b111011101110;
20'b01000110100011011000: color_data = 12'b111011101110;
20'b01000110100011011001: color_data = 12'b111011101110;
20'b01000110100011011010: color_data = 12'b111011101110;
20'b01000110100011011011: color_data = 12'b111011101110;
20'b01000110100011011100: color_data = 12'b111011101110;
20'b01000110100011011101: color_data = 12'b111011101110;
20'b01000110100011011110: color_data = 12'b111011101110;
20'b01000110100011011111: color_data = 12'b111011101110;
20'b01000110100011100000: color_data = 12'b111011101110;
20'b01000110100011100001: color_data = 12'b111011101110;
20'b01000110100011101101: color_data = 12'b111011101110;
20'b01000110100011101110: color_data = 12'b111011101110;
20'b01000110100011101111: color_data = 12'b111011101110;
20'b01000110100011110000: color_data = 12'b111011101110;
20'b01000110100011110001: color_data = 12'b111011101110;
20'b01000110100011110010: color_data = 12'b111011101110;
20'b01000110100011110011: color_data = 12'b111011101110;
20'b01000110100011110100: color_data = 12'b111011101110;
20'b01000110100011110101: color_data = 12'b111011101110;
20'b01000110100011110110: color_data = 12'b111011101110;
20'b01000110100011111000: color_data = 12'b111011101110;
20'b01000110100011111001: color_data = 12'b111011101110;
20'b01000110100011111010: color_data = 12'b111011101110;
20'b01000110100011111011: color_data = 12'b111011101110;
20'b01000110100011111100: color_data = 12'b111011101110;
20'b01000110100011111101: color_data = 12'b111011101110;
20'b01000110100011111110: color_data = 12'b111011101110;
20'b01000110100011111111: color_data = 12'b111011101110;
20'b01000110100100000000: color_data = 12'b111011101110;
20'b01000110100100000001: color_data = 12'b111011101110;
20'b01000110100100100100: color_data = 12'b111011101110;
20'b01000110100100100101: color_data = 12'b111011101110;
20'b01000110100100100110: color_data = 12'b111011101110;
20'b01000110100100100111: color_data = 12'b111011101110;
20'b01000110100100101000: color_data = 12'b111011101110;
20'b01000110100100101001: color_data = 12'b111011101110;
20'b01000110100100101010: color_data = 12'b111011101110;
20'b01000110100100101011: color_data = 12'b111011101110;
20'b01000110100100101100: color_data = 12'b111011101110;
20'b01000110100100101101: color_data = 12'b111011101110;
20'b01000110100100101111: color_data = 12'b111011101110;
20'b01000110100100110000: color_data = 12'b111011101110;
20'b01000110100100110001: color_data = 12'b111011101110;
20'b01000110100100110010: color_data = 12'b111011101110;
20'b01000110100100110011: color_data = 12'b111011101110;
20'b01000110100100110100: color_data = 12'b111011101110;
20'b01000110100100110101: color_data = 12'b111011101110;
20'b01000110100100110110: color_data = 12'b111011101110;
20'b01000110100100110111: color_data = 12'b111011101110;
20'b01000110100100111000: color_data = 12'b111011101110;
20'b01000110100101000100: color_data = 12'b111011101110;
20'b01000110100101000101: color_data = 12'b111011101110;
20'b01000110100101000110: color_data = 12'b111011101110;
20'b01000110100101000111: color_data = 12'b111011101110;
20'b01000110100101001000: color_data = 12'b111011101110;
20'b01000110100101001001: color_data = 12'b111011101110;
20'b01000110100101001010: color_data = 12'b111011101110;
20'b01000110100101001011: color_data = 12'b111011101110;
20'b01000110100101001100: color_data = 12'b111011101110;
20'b01000110100101001101: color_data = 12'b111011101110;
20'b01000110100101001111: color_data = 12'b111011101110;
20'b01000110100101010000: color_data = 12'b111011101110;
20'b01000110100101010001: color_data = 12'b111011101110;
20'b01000110100101010010: color_data = 12'b111011101110;
20'b01000110100101010011: color_data = 12'b111011101110;
20'b01000110100101010100: color_data = 12'b111011101110;
20'b01000110100101010101: color_data = 12'b111011101110;
20'b01000110100101010110: color_data = 12'b111011101110;
20'b01000110100101010111: color_data = 12'b111011101110;
20'b01000110100101011000: color_data = 12'b111011101110;
20'b01000110100110011100: color_data = 12'b111011101110;
20'b01000110100110011101: color_data = 12'b111011101110;
20'b01000110100110011110: color_data = 12'b111011101110;
20'b01000110100110011111: color_data = 12'b111011101110;
20'b01000110100110100000: color_data = 12'b111011101110;
20'b01000110100110100001: color_data = 12'b111011101110;
20'b01000110100110100010: color_data = 12'b111011101110;
20'b01000110100110100011: color_data = 12'b111011101110;
20'b01000110100110100100: color_data = 12'b111011101110;
20'b01000110100110100101: color_data = 12'b111011101110;
20'b01000110100110100111: color_data = 12'b111011101110;
20'b01000110100110101000: color_data = 12'b111011101110;
20'b01000110100110101001: color_data = 12'b111011101110;
20'b01000110100110101010: color_data = 12'b111011101110;
20'b01000110100110101011: color_data = 12'b111011101110;
20'b01000110100110101100: color_data = 12'b111011101110;
20'b01000110100110101101: color_data = 12'b111011101110;
20'b01000110100110101110: color_data = 12'b111011101110;
20'b01000110100110101111: color_data = 12'b111011101110;
20'b01000110100110110000: color_data = 12'b111011101110;
20'b01000110100111010011: color_data = 12'b111011101110;
20'b01000110100111010100: color_data = 12'b111011101110;
20'b01000110100111010101: color_data = 12'b111011101110;
20'b01000110100111010110: color_data = 12'b111011101110;
20'b01000110100111010111: color_data = 12'b111011101110;
20'b01000110100111011000: color_data = 12'b111011101110;
20'b01000110100111011001: color_data = 12'b111011101110;
20'b01000110100111011010: color_data = 12'b111011101110;
20'b01000110100111011011: color_data = 12'b111011101110;
20'b01000110100111011100: color_data = 12'b111011101110;
20'b01000110100111011110: color_data = 12'b111011101110;
20'b01000110100111011111: color_data = 12'b111011101110;
20'b01000110100111100000: color_data = 12'b111011101110;
20'b01000110100111100001: color_data = 12'b111011101110;
20'b01000110100111100010: color_data = 12'b111011101110;
20'b01000110100111100011: color_data = 12'b111011101110;
20'b01000110100111100100: color_data = 12'b111011101110;
20'b01000110100111100101: color_data = 12'b111011101110;
20'b01000110100111100110: color_data = 12'b111011101110;
20'b01000110100111100111: color_data = 12'b111011101110;
20'b01000110110010010110: color_data = 12'b111011101110;
20'b01000110110010010111: color_data = 12'b111011101110;
20'b01000110110010011000: color_data = 12'b111011101110;
20'b01000110110010011001: color_data = 12'b111011101110;
20'b01000110110010011010: color_data = 12'b111011101110;
20'b01000110110010011011: color_data = 12'b111011101110;
20'b01000110110010011100: color_data = 12'b111011101110;
20'b01000110110010011101: color_data = 12'b111011101110;
20'b01000110110010011110: color_data = 12'b111011101110;
20'b01000110110010011111: color_data = 12'b111011101110;
20'b01000110110010100001: color_data = 12'b111011101110;
20'b01000110110010100010: color_data = 12'b111011101110;
20'b01000110110010100011: color_data = 12'b111011101110;
20'b01000110110010100100: color_data = 12'b111011101110;
20'b01000110110010100101: color_data = 12'b111011101110;
20'b01000110110010100110: color_data = 12'b111011101110;
20'b01000110110010100111: color_data = 12'b111011101110;
20'b01000110110010101000: color_data = 12'b111011101110;
20'b01000110110010101001: color_data = 12'b111011101110;
20'b01000110110010101010: color_data = 12'b111011101110;
20'b01000110110011001101: color_data = 12'b111011101110;
20'b01000110110011001110: color_data = 12'b111011101110;
20'b01000110110011001111: color_data = 12'b111011101110;
20'b01000110110011010000: color_data = 12'b111011101110;
20'b01000110110011010001: color_data = 12'b111011101110;
20'b01000110110011010010: color_data = 12'b111011101110;
20'b01000110110011010011: color_data = 12'b111011101110;
20'b01000110110011010100: color_data = 12'b111011101110;
20'b01000110110011010101: color_data = 12'b111011101110;
20'b01000110110011010110: color_data = 12'b111011101110;
20'b01000110110011011000: color_data = 12'b111011101110;
20'b01000110110011011001: color_data = 12'b111011101110;
20'b01000110110011011010: color_data = 12'b111011101110;
20'b01000110110011011011: color_data = 12'b111011101110;
20'b01000110110011011100: color_data = 12'b111011101110;
20'b01000110110011011101: color_data = 12'b111011101110;
20'b01000110110011011110: color_data = 12'b111011101110;
20'b01000110110011011111: color_data = 12'b111011101110;
20'b01000110110011100000: color_data = 12'b111011101110;
20'b01000110110011100001: color_data = 12'b111011101110;
20'b01000110110011101101: color_data = 12'b111011101110;
20'b01000110110011101110: color_data = 12'b111011101110;
20'b01000110110011101111: color_data = 12'b111011101110;
20'b01000110110011110000: color_data = 12'b111011101110;
20'b01000110110011110001: color_data = 12'b111011101110;
20'b01000110110011110010: color_data = 12'b111011101110;
20'b01000110110011110011: color_data = 12'b111011101110;
20'b01000110110011110100: color_data = 12'b111011101110;
20'b01000110110011110101: color_data = 12'b111011101110;
20'b01000110110011110110: color_data = 12'b111011101110;
20'b01000110110011111000: color_data = 12'b111011101110;
20'b01000110110011111001: color_data = 12'b111011101110;
20'b01000110110011111010: color_data = 12'b111011101110;
20'b01000110110011111011: color_data = 12'b111011101110;
20'b01000110110011111100: color_data = 12'b111011101110;
20'b01000110110011111101: color_data = 12'b111011101110;
20'b01000110110011111110: color_data = 12'b111011101110;
20'b01000110110011111111: color_data = 12'b111011101110;
20'b01000110110100000000: color_data = 12'b111011101110;
20'b01000110110100000001: color_data = 12'b111011101110;
20'b01000110110100100100: color_data = 12'b111011101110;
20'b01000110110100100101: color_data = 12'b111011101110;
20'b01000110110100100110: color_data = 12'b111011101110;
20'b01000110110100100111: color_data = 12'b111011101110;
20'b01000110110100101000: color_data = 12'b111011101110;
20'b01000110110100101001: color_data = 12'b111011101110;
20'b01000110110100101010: color_data = 12'b111011101110;
20'b01000110110100101011: color_data = 12'b111011101110;
20'b01000110110100101100: color_data = 12'b111011101110;
20'b01000110110100101101: color_data = 12'b111011101110;
20'b01000110110100101111: color_data = 12'b111011101110;
20'b01000110110100110000: color_data = 12'b111011101110;
20'b01000110110100110001: color_data = 12'b111011101110;
20'b01000110110100110010: color_data = 12'b111011101110;
20'b01000110110100110011: color_data = 12'b111011101110;
20'b01000110110100110100: color_data = 12'b111011101110;
20'b01000110110100110101: color_data = 12'b111011101110;
20'b01000110110100110110: color_data = 12'b111011101110;
20'b01000110110100110111: color_data = 12'b111011101110;
20'b01000110110100111000: color_data = 12'b111011101110;
20'b01000110110101000100: color_data = 12'b111011101110;
20'b01000110110101000101: color_data = 12'b111011101110;
20'b01000110110101000110: color_data = 12'b111011101110;
20'b01000110110101000111: color_data = 12'b111011101110;
20'b01000110110101001000: color_data = 12'b111011101110;
20'b01000110110101001001: color_data = 12'b111011101110;
20'b01000110110101001010: color_data = 12'b111011101110;
20'b01000110110101001011: color_data = 12'b111011101110;
20'b01000110110101001100: color_data = 12'b111011101110;
20'b01000110110101001101: color_data = 12'b111011101110;
20'b01000110110101001111: color_data = 12'b111011101110;
20'b01000110110101010000: color_data = 12'b111011101110;
20'b01000110110101010001: color_data = 12'b111011101110;
20'b01000110110101010010: color_data = 12'b111011101110;
20'b01000110110101010011: color_data = 12'b111011101110;
20'b01000110110101010100: color_data = 12'b111011101110;
20'b01000110110101010101: color_data = 12'b111011101110;
20'b01000110110101010110: color_data = 12'b111011101110;
20'b01000110110101010111: color_data = 12'b111011101110;
20'b01000110110101011000: color_data = 12'b111011101110;
20'b01000110110110011100: color_data = 12'b111011101110;
20'b01000110110110011101: color_data = 12'b111011101110;
20'b01000110110110011110: color_data = 12'b111011101110;
20'b01000110110110011111: color_data = 12'b111011101110;
20'b01000110110110100000: color_data = 12'b111011101110;
20'b01000110110110100001: color_data = 12'b111011101110;
20'b01000110110110100010: color_data = 12'b111011101110;
20'b01000110110110100011: color_data = 12'b111011101110;
20'b01000110110110100100: color_data = 12'b111011101110;
20'b01000110110110100101: color_data = 12'b111011101110;
20'b01000110110110100111: color_data = 12'b111011101110;
20'b01000110110110101000: color_data = 12'b111011101110;
20'b01000110110110101001: color_data = 12'b111011101110;
20'b01000110110110101010: color_data = 12'b111011101110;
20'b01000110110110101011: color_data = 12'b111011101110;
20'b01000110110110101100: color_data = 12'b111011101110;
20'b01000110110110101101: color_data = 12'b111011101110;
20'b01000110110110101110: color_data = 12'b111011101110;
20'b01000110110110101111: color_data = 12'b111011101110;
20'b01000110110110110000: color_data = 12'b111011101110;
20'b01000110110111010011: color_data = 12'b111011101110;
20'b01000110110111010100: color_data = 12'b111011101110;
20'b01000110110111010101: color_data = 12'b111011101110;
20'b01000110110111010110: color_data = 12'b111011101110;
20'b01000110110111010111: color_data = 12'b111011101110;
20'b01000110110111011000: color_data = 12'b111011101110;
20'b01000110110111011001: color_data = 12'b111011101110;
20'b01000110110111011010: color_data = 12'b111011101110;
20'b01000110110111011011: color_data = 12'b111011101110;
20'b01000110110111011100: color_data = 12'b111011101110;
20'b01000110110111011110: color_data = 12'b111011101110;
20'b01000110110111011111: color_data = 12'b111011101110;
20'b01000110110111100000: color_data = 12'b111011101110;
20'b01000110110111100001: color_data = 12'b111011101110;
20'b01000110110111100010: color_data = 12'b111011101110;
20'b01000110110111100011: color_data = 12'b111011101110;
20'b01000110110111100100: color_data = 12'b111011101110;
20'b01000110110111100101: color_data = 12'b111011101110;
20'b01000110110111100110: color_data = 12'b111011101110;
20'b01000110110111100111: color_data = 12'b111011101110;
20'b01000111000010010110: color_data = 12'b111011101110;
20'b01000111000010010111: color_data = 12'b111011101110;
20'b01000111000010011000: color_data = 12'b111011101110;
20'b01000111000010011001: color_data = 12'b111011101110;
20'b01000111000010011010: color_data = 12'b111011101110;
20'b01000111000010011011: color_data = 12'b111011101110;
20'b01000111000010011100: color_data = 12'b111011101110;
20'b01000111000010011101: color_data = 12'b111011101110;
20'b01000111000010011110: color_data = 12'b111011101110;
20'b01000111000010011111: color_data = 12'b111011101110;
20'b01000111000010100001: color_data = 12'b111011101110;
20'b01000111000010100010: color_data = 12'b111011101110;
20'b01000111000010100011: color_data = 12'b111011101110;
20'b01000111000010100100: color_data = 12'b111011101110;
20'b01000111000010100101: color_data = 12'b111011101110;
20'b01000111000010100110: color_data = 12'b111011101110;
20'b01000111000010100111: color_data = 12'b111011101110;
20'b01000111000010101000: color_data = 12'b111011101110;
20'b01000111000010101001: color_data = 12'b111011101110;
20'b01000111000010101010: color_data = 12'b111011101110;
20'b01000111000011001101: color_data = 12'b111011101110;
20'b01000111000011001110: color_data = 12'b111011101110;
20'b01000111000011001111: color_data = 12'b111011101110;
20'b01000111000011010000: color_data = 12'b111011101110;
20'b01000111000011010001: color_data = 12'b111011101110;
20'b01000111000011010010: color_data = 12'b111011101110;
20'b01000111000011010011: color_data = 12'b111011101110;
20'b01000111000011010100: color_data = 12'b111011101110;
20'b01000111000011010101: color_data = 12'b111011101110;
20'b01000111000011010110: color_data = 12'b111011101110;
20'b01000111000011011000: color_data = 12'b111011101110;
20'b01000111000011011001: color_data = 12'b111011101110;
20'b01000111000011011010: color_data = 12'b111011101110;
20'b01000111000011011011: color_data = 12'b111011101110;
20'b01000111000011011100: color_data = 12'b111011101110;
20'b01000111000011011101: color_data = 12'b111011101110;
20'b01000111000011011110: color_data = 12'b111011101110;
20'b01000111000011011111: color_data = 12'b111011101110;
20'b01000111000011100000: color_data = 12'b111011101110;
20'b01000111000011100001: color_data = 12'b111011101110;
20'b01000111000011101101: color_data = 12'b111011101110;
20'b01000111000011101110: color_data = 12'b111011101110;
20'b01000111000011101111: color_data = 12'b111011101110;
20'b01000111000011110000: color_data = 12'b111011101110;
20'b01000111000011110001: color_data = 12'b111011101110;
20'b01000111000011110010: color_data = 12'b111011101110;
20'b01000111000011110011: color_data = 12'b111011101110;
20'b01000111000011110100: color_data = 12'b111011101110;
20'b01000111000011110101: color_data = 12'b111011101110;
20'b01000111000011110110: color_data = 12'b111011101110;
20'b01000111000011111000: color_data = 12'b111011101110;
20'b01000111000011111001: color_data = 12'b111011101110;
20'b01000111000011111010: color_data = 12'b111011101110;
20'b01000111000011111011: color_data = 12'b111011101110;
20'b01000111000011111100: color_data = 12'b111011101110;
20'b01000111000011111101: color_data = 12'b111011101110;
20'b01000111000011111110: color_data = 12'b111011101110;
20'b01000111000011111111: color_data = 12'b111011101110;
20'b01000111000100000000: color_data = 12'b111011101110;
20'b01000111000100000001: color_data = 12'b111011101110;
20'b01000111000100100100: color_data = 12'b111011101110;
20'b01000111000100100101: color_data = 12'b111011101110;
20'b01000111000100100110: color_data = 12'b111011101110;
20'b01000111000100100111: color_data = 12'b111011101110;
20'b01000111000100101000: color_data = 12'b111011101110;
20'b01000111000100101001: color_data = 12'b111011101110;
20'b01000111000100101010: color_data = 12'b111011101110;
20'b01000111000100101011: color_data = 12'b111011101110;
20'b01000111000100101100: color_data = 12'b111011101110;
20'b01000111000100101101: color_data = 12'b111011101110;
20'b01000111000100101111: color_data = 12'b111011101110;
20'b01000111000100110000: color_data = 12'b111011101110;
20'b01000111000100110001: color_data = 12'b111011101110;
20'b01000111000100110010: color_data = 12'b111011101110;
20'b01000111000100110011: color_data = 12'b111011101110;
20'b01000111000100110100: color_data = 12'b111011101110;
20'b01000111000100110101: color_data = 12'b111011101110;
20'b01000111000100110110: color_data = 12'b111011101110;
20'b01000111000100110111: color_data = 12'b111011101110;
20'b01000111000100111000: color_data = 12'b111011101110;
20'b01000111000101000100: color_data = 12'b111011101110;
20'b01000111000101000101: color_data = 12'b111011101110;
20'b01000111000101000110: color_data = 12'b111011101110;
20'b01000111000101000111: color_data = 12'b111011101110;
20'b01000111000101001000: color_data = 12'b111011101110;
20'b01000111000101001001: color_data = 12'b111011101110;
20'b01000111000101001010: color_data = 12'b111011101110;
20'b01000111000101001011: color_data = 12'b111011101110;
20'b01000111000101001100: color_data = 12'b111011101110;
20'b01000111000101001101: color_data = 12'b111011101110;
20'b01000111000101001111: color_data = 12'b111011101110;
20'b01000111000101010000: color_data = 12'b111011101110;
20'b01000111000101010001: color_data = 12'b111011101110;
20'b01000111000101010010: color_data = 12'b111011101110;
20'b01000111000101010011: color_data = 12'b111011101110;
20'b01000111000101010100: color_data = 12'b111011101110;
20'b01000111000101010101: color_data = 12'b111011101110;
20'b01000111000101010110: color_data = 12'b111011101110;
20'b01000111000101010111: color_data = 12'b111011101110;
20'b01000111000101011000: color_data = 12'b111011101110;
20'b01000111000110011100: color_data = 12'b111011101110;
20'b01000111000110011101: color_data = 12'b111011101110;
20'b01000111000110011110: color_data = 12'b111011101110;
20'b01000111000110011111: color_data = 12'b111011101110;
20'b01000111000110100000: color_data = 12'b111011101110;
20'b01000111000110100001: color_data = 12'b111011101110;
20'b01000111000110100010: color_data = 12'b111011101110;
20'b01000111000110100011: color_data = 12'b111011101110;
20'b01000111000110100100: color_data = 12'b111011101110;
20'b01000111000110100101: color_data = 12'b111011101110;
20'b01000111000110100111: color_data = 12'b111011101110;
20'b01000111000110101000: color_data = 12'b111011101110;
20'b01000111000110101001: color_data = 12'b111011101110;
20'b01000111000110101010: color_data = 12'b111011101110;
20'b01000111000110101011: color_data = 12'b111011101110;
20'b01000111000110101100: color_data = 12'b111011101110;
20'b01000111000110101101: color_data = 12'b111011101110;
20'b01000111000110101110: color_data = 12'b111011101110;
20'b01000111000110101111: color_data = 12'b111011101110;
20'b01000111000110110000: color_data = 12'b111011101110;
20'b01000111000111010011: color_data = 12'b111011101110;
20'b01000111000111010100: color_data = 12'b111011101110;
20'b01000111000111010101: color_data = 12'b111011101110;
20'b01000111000111010110: color_data = 12'b111011101110;
20'b01000111000111010111: color_data = 12'b111011101110;
20'b01000111000111011000: color_data = 12'b111011101110;
20'b01000111000111011001: color_data = 12'b111011101110;
20'b01000111000111011010: color_data = 12'b111011101110;
20'b01000111000111011011: color_data = 12'b111011101110;
20'b01000111000111011100: color_data = 12'b111011101110;
20'b01000111000111011110: color_data = 12'b111011101110;
20'b01000111000111011111: color_data = 12'b111011101110;
20'b01000111000111100000: color_data = 12'b111011101110;
20'b01000111000111100001: color_data = 12'b111011101110;
20'b01000111000111100010: color_data = 12'b111011101110;
20'b01000111000111100011: color_data = 12'b111011101110;
20'b01000111000111100100: color_data = 12'b111011101110;
20'b01000111000111100101: color_data = 12'b111011101110;
20'b01000111000111100110: color_data = 12'b111011101110;
20'b01000111000111100111: color_data = 12'b111011101110;
20'b01000111010010010110: color_data = 12'b111011101110;
20'b01000111010010010111: color_data = 12'b111011101110;
20'b01000111010010011000: color_data = 12'b111011101110;
20'b01000111010010011001: color_data = 12'b111011101110;
20'b01000111010010011010: color_data = 12'b111011101110;
20'b01000111010010011011: color_data = 12'b111011101110;
20'b01000111010010011100: color_data = 12'b111011101110;
20'b01000111010010011101: color_data = 12'b111011101110;
20'b01000111010010011110: color_data = 12'b111011101110;
20'b01000111010010011111: color_data = 12'b111011101110;
20'b01000111010010100001: color_data = 12'b111011101110;
20'b01000111010010100010: color_data = 12'b111011101110;
20'b01000111010010100011: color_data = 12'b111011101110;
20'b01000111010010100100: color_data = 12'b111011101110;
20'b01000111010010100101: color_data = 12'b111011101110;
20'b01000111010010100110: color_data = 12'b111011101110;
20'b01000111010010100111: color_data = 12'b111011101110;
20'b01000111010010101000: color_data = 12'b111011101110;
20'b01000111010010101001: color_data = 12'b111011101110;
20'b01000111010010101010: color_data = 12'b111011101110;
20'b01000111010011001101: color_data = 12'b111011101110;
20'b01000111010011001110: color_data = 12'b111011101110;
20'b01000111010011001111: color_data = 12'b111011101110;
20'b01000111010011010000: color_data = 12'b111011101110;
20'b01000111010011010001: color_data = 12'b111011101110;
20'b01000111010011010010: color_data = 12'b111011101110;
20'b01000111010011010011: color_data = 12'b111011101110;
20'b01000111010011010100: color_data = 12'b111011101110;
20'b01000111010011010101: color_data = 12'b111011101110;
20'b01000111010011010110: color_data = 12'b111011101110;
20'b01000111010011011000: color_data = 12'b111011101110;
20'b01000111010011011001: color_data = 12'b111011101110;
20'b01000111010011011010: color_data = 12'b111011101110;
20'b01000111010011011011: color_data = 12'b111011101110;
20'b01000111010011011100: color_data = 12'b111011101110;
20'b01000111010011011101: color_data = 12'b111011101110;
20'b01000111010011011110: color_data = 12'b111011101110;
20'b01000111010011011111: color_data = 12'b111011101110;
20'b01000111010011100000: color_data = 12'b111011101110;
20'b01000111010011100001: color_data = 12'b111011101110;
20'b01000111010011101101: color_data = 12'b111011101110;
20'b01000111010011101110: color_data = 12'b111011101110;
20'b01000111010011101111: color_data = 12'b111011101110;
20'b01000111010011110000: color_data = 12'b111011101110;
20'b01000111010011110001: color_data = 12'b111011101110;
20'b01000111010011110010: color_data = 12'b111011101110;
20'b01000111010011110011: color_data = 12'b111011101110;
20'b01000111010011110100: color_data = 12'b111011101110;
20'b01000111010011110101: color_data = 12'b111011101110;
20'b01000111010011110110: color_data = 12'b111011101110;
20'b01000111010011111000: color_data = 12'b111011101110;
20'b01000111010011111001: color_data = 12'b111011101110;
20'b01000111010011111010: color_data = 12'b111011101110;
20'b01000111010011111011: color_data = 12'b111011101110;
20'b01000111010011111100: color_data = 12'b111011101110;
20'b01000111010011111101: color_data = 12'b111011101110;
20'b01000111010011111110: color_data = 12'b111011101110;
20'b01000111010011111111: color_data = 12'b111011101110;
20'b01000111010100000000: color_data = 12'b111011101110;
20'b01000111010100000001: color_data = 12'b111011101110;
20'b01000111010100100100: color_data = 12'b111011101110;
20'b01000111010100100101: color_data = 12'b111011101110;
20'b01000111010100100110: color_data = 12'b111011101110;
20'b01000111010100100111: color_data = 12'b111011101110;
20'b01000111010100101000: color_data = 12'b111011101110;
20'b01000111010100101001: color_data = 12'b111011101110;
20'b01000111010100101010: color_data = 12'b111011101110;
20'b01000111010100101011: color_data = 12'b111011101110;
20'b01000111010100101100: color_data = 12'b111011101110;
20'b01000111010100101101: color_data = 12'b111011101110;
20'b01000111010100101111: color_data = 12'b111011101110;
20'b01000111010100110000: color_data = 12'b111011101110;
20'b01000111010100110001: color_data = 12'b111011101110;
20'b01000111010100110010: color_data = 12'b111011101110;
20'b01000111010100110011: color_data = 12'b111011101110;
20'b01000111010100110100: color_data = 12'b111011101110;
20'b01000111010100110101: color_data = 12'b111011101110;
20'b01000111010100110110: color_data = 12'b111011101110;
20'b01000111010100110111: color_data = 12'b111011101110;
20'b01000111010100111000: color_data = 12'b111011101110;
20'b01000111010101000100: color_data = 12'b111011101110;
20'b01000111010101000101: color_data = 12'b111011101110;
20'b01000111010101000110: color_data = 12'b111011101110;
20'b01000111010101000111: color_data = 12'b111011101110;
20'b01000111010101001000: color_data = 12'b111011101110;
20'b01000111010101001001: color_data = 12'b111011101110;
20'b01000111010101001010: color_data = 12'b111011101110;
20'b01000111010101001011: color_data = 12'b111011101110;
20'b01000111010101001100: color_data = 12'b111011101110;
20'b01000111010101001101: color_data = 12'b111011101110;
20'b01000111010101001111: color_data = 12'b111011101110;
20'b01000111010101010000: color_data = 12'b111011101110;
20'b01000111010101010001: color_data = 12'b111011101110;
20'b01000111010101010010: color_data = 12'b111011101110;
20'b01000111010101010011: color_data = 12'b111011101110;
20'b01000111010101010100: color_data = 12'b111011101110;
20'b01000111010101010101: color_data = 12'b111011101110;
20'b01000111010101010110: color_data = 12'b111011101110;
20'b01000111010101010111: color_data = 12'b111011101110;
20'b01000111010101011000: color_data = 12'b111011101110;
20'b01000111010110011100: color_data = 12'b111011101110;
20'b01000111010110011101: color_data = 12'b111011101110;
20'b01000111010110011110: color_data = 12'b111011101110;
20'b01000111010110011111: color_data = 12'b111011101110;
20'b01000111010110100000: color_data = 12'b111011101110;
20'b01000111010110100001: color_data = 12'b111011101110;
20'b01000111010110100010: color_data = 12'b111011101110;
20'b01000111010110100011: color_data = 12'b111011101110;
20'b01000111010110100100: color_data = 12'b111011101110;
20'b01000111010110100101: color_data = 12'b111011101110;
20'b01000111010110100111: color_data = 12'b111011101110;
20'b01000111010110101000: color_data = 12'b111011101110;
20'b01000111010110101001: color_data = 12'b111011101110;
20'b01000111010110101010: color_data = 12'b111011101110;
20'b01000111010110101011: color_data = 12'b111011101110;
20'b01000111010110101100: color_data = 12'b111011101110;
20'b01000111010110101101: color_data = 12'b111011101110;
20'b01000111010110101110: color_data = 12'b111011101110;
20'b01000111010110101111: color_data = 12'b111011101110;
20'b01000111010110110000: color_data = 12'b111011101110;
20'b01000111010111010011: color_data = 12'b111011101110;
20'b01000111010111010100: color_data = 12'b111011101110;
20'b01000111010111010101: color_data = 12'b111011101110;
20'b01000111010111010110: color_data = 12'b111011101110;
20'b01000111010111010111: color_data = 12'b111011101110;
20'b01000111010111011000: color_data = 12'b111011101110;
20'b01000111010111011001: color_data = 12'b111011101110;
20'b01000111010111011010: color_data = 12'b111011101110;
20'b01000111010111011011: color_data = 12'b111011101110;
20'b01000111010111011100: color_data = 12'b111011101110;
20'b01000111010111011110: color_data = 12'b111011101110;
20'b01000111010111011111: color_data = 12'b111011101110;
20'b01000111010111100000: color_data = 12'b111011101110;
20'b01000111010111100001: color_data = 12'b111011101110;
20'b01000111010111100010: color_data = 12'b111011101110;
20'b01000111010111100011: color_data = 12'b111011101110;
20'b01000111010111100100: color_data = 12'b111011101110;
20'b01000111010111100101: color_data = 12'b111011101110;
20'b01000111010111100110: color_data = 12'b111011101110;
20'b01000111010111100111: color_data = 12'b111011101110;
20'b01000111100010010110: color_data = 12'b111011101110;
20'b01000111100010010111: color_data = 12'b111011101110;
20'b01000111100010011000: color_data = 12'b111011101110;
20'b01000111100010011001: color_data = 12'b111011101110;
20'b01000111100010011010: color_data = 12'b111011101110;
20'b01000111100010011011: color_data = 12'b111011101110;
20'b01000111100010011100: color_data = 12'b111011101110;
20'b01000111100010011101: color_data = 12'b111011101110;
20'b01000111100010011110: color_data = 12'b111011101110;
20'b01000111100010011111: color_data = 12'b111011101110;
20'b01000111100010100001: color_data = 12'b111011101110;
20'b01000111100010100010: color_data = 12'b111011101110;
20'b01000111100010100011: color_data = 12'b111011101110;
20'b01000111100010100100: color_data = 12'b111011101110;
20'b01000111100010100101: color_data = 12'b111011101110;
20'b01000111100010100110: color_data = 12'b111011101110;
20'b01000111100010100111: color_data = 12'b111011101110;
20'b01000111100010101000: color_data = 12'b111011101110;
20'b01000111100010101001: color_data = 12'b111011101110;
20'b01000111100010101010: color_data = 12'b111011101110;
20'b01000111100011001101: color_data = 12'b111011101110;
20'b01000111100011001110: color_data = 12'b111011101110;
20'b01000111100011001111: color_data = 12'b111011101110;
20'b01000111100011010000: color_data = 12'b111011101110;
20'b01000111100011010001: color_data = 12'b111011101110;
20'b01000111100011010010: color_data = 12'b111011101110;
20'b01000111100011010011: color_data = 12'b111011101110;
20'b01000111100011010100: color_data = 12'b111011101110;
20'b01000111100011010101: color_data = 12'b111011101110;
20'b01000111100011010110: color_data = 12'b111011101110;
20'b01000111100011011000: color_data = 12'b111011101110;
20'b01000111100011011001: color_data = 12'b111011101110;
20'b01000111100011011010: color_data = 12'b111011101110;
20'b01000111100011011011: color_data = 12'b111011101110;
20'b01000111100011011100: color_data = 12'b111011101110;
20'b01000111100011011101: color_data = 12'b111011101110;
20'b01000111100011011110: color_data = 12'b111011101110;
20'b01000111100011011111: color_data = 12'b111011101110;
20'b01000111100011100000: color_data = 12'b111011101110;
20'b01000111100011100001: color_data = 12'b111011101110;
20'b01000111100011101101: color_data = 12'b111011101110;
20'b01000111100011101110: color_data = 12'b111011101110;
20'b01000111100011101111: color_data = 12'b111011101110;
20'b01000111100011110000: color_data = 12'b111011101110;
20'b01000111100011110001: color_data = 12'b111011101110;
20'b01000111100011110010: color_data = 12'b111011101110;
20'b01000111100011110011: color_data = 12'b111011101110;
20'b01000111100011110100: color_data = 12'b111011101110;
20'b01000111100011110101: color_data = 12'b111011101110;
20'b01000111100011110110: color_data = 12'b111011101110;
20'b01000111100011111000: color_data = 12'b111011101110;
20'b01000111100011111001: color_data = 12'b111011101110;
20'b01000111100011111010: color_data = 12'b111011101110;
20'b01000111100011111011: color_data = 12'b111011101110;
20'b01000111100011111100: color_data = 12'b111011101110;
20'b01000111100011111101: color_data = 12'b111011101110;
20'b01000111100011111110: color_data = 12'b111011101110;
20'b01000111100011111111: color_data = 12'b111011101110;
20'b01000111100100000000: color_data = 12'b111011101110;
20'b01000111100100000001: color_data = 12'b111011101110;
20'b01000111100100100100: color_data = 12'b111011101110;
20'b01000111100100100101: color_data = 12'b111011101110;
20'b01000111100100100110: color_data = 12'b111011101110;
20'b01000111100100100111: color_data = 12'b111011101110;
20'b01000111100100101000: color_data = 12'b111011101110;
20'b01000111100100101001: color_data = 12'b111011101110;
20'b01000111100100101010: color_data = 12'b111011101110;
20'b01000111100100101011: color_data = 12'b111011101110;
20'b01000111100100101100: color_data = 12'b111011101110;
20'b01000111100100101101: color_data = 12'b111011101110;
20'b01000111100100101111: color_data = 12'b111011101110;
20'b01000111100100110000: color_data = 12'b111011101110;
20'b01000111100100110001: color_data = 12'b111011101110;
20'b01000111100100110010: color_data = 12'b111011101110;
20'b01000111100100110011: color_data = 12'b111011101110;
20'b01000111100100110100: color_data = 12'b111011101110;
20'b01000111100100110101: color_data = 12'b111011101110;
20'b01000111100100110110: color_data = 12'b111011101110;
20'b01000111100100110111: color_data = 12'b111011101110;
20'b01000111100100111000: color_data = 12'b111011101110;
20'b01000111100101000100: color_data = 12'b111011101110;
20'b01000111100101000101: color_data = 12'b111011101110;
20'b01000111100101000110: color_data = 12'b111011101110;
20'b01000111100101000111: color_data = 12'b111011101110;
20'b01000111100101001000: color_data = 12'b111011101110;
20'b01000111100101001001: color_data = 12'b111011101110;
20'b01000111100101001010: color_data = 12'b111011101110;
20'b01000111100101001011: color_data = 12'b111011101110;
20'b01000111100101001100: color_data = 12'b111011101110;
20'b01000111100101001101: color_data = 12'b111011101110;
20'b01000111100101001111: color_data = 12'b111011101110;
20'b01000111100101010000: color_data = 12'b111011101110;
20'b01000111100101010001: color_data = 12'b111011101110;
20'b01000111100101010010: color_data = 12'b111011101110;
20'b01000111100101010011: color_data = 12'b111011101110;
20'b01000111100101010100: color_data = 12'b111011101110;
20'b01000111100101010101: color_data = 12'b111011101110;
20'b01000111100101010110: color_data = 12'b111011101110;
20'b01000111100101010111: color_data = 12'b111011101110;
20'b01000111100101011000: color_data = 12'b111011101110;
20'b01000111100110011100: color_data = 12'b111011101110;
20'b01000111100110011101: color_data = 12'b111011101110;
20'b01000111100110011110: color_data = 12'b111011101110;
20'b01000111100110011111: color_data = 12'b111011101110;
20'b01000111100110100000: color_data = 12'b111011101110;
20'b01000111100110100001: color_data = 12'b111011101110;
20'b01000111100110100010: color_data = 12'b111011101110;
20'b01000111100110100011: color_data = 12'b111011101110;
20'b01000111100110100100: color_data = 12'b111011101110;
20'b01000111100110100101: color_data = 12'b111011101110;
20'b01000111100110100111: color_data = 12'b111011101110;
20'b01000111100110101000: color_data = 12'b111011101110;
20'b01000111100110101001: color_data = 12'b111011101110;
20'b01000111100110101010: color_data = 12'b111011101110;
20'b01000111100110101011: color_data = 12'b111011101110;
20'b01000111100110101100: color_data = 12'b111011101110;
20'b01000111100110101101: color_data = 12'b111011101110;
20'b01000111100110101110: color_data = 12'b111011101110;
20'b01000111100110101111: color_data = 12'b111011101110;
20'b01000111100110110000: color_data = 12'b111011101110;
20'b01000111100111010011: color_data = 12'b111011101110;
20'b01000111100111010100: color_data = 12'b111011101110;
20'b01000111100111010101: color_data = 12'b111011101110;
20'b01000111100111010110: color_data = 12'b111011101110;
20'b01000111100111010111: color_data = 12'b111011101110;
20'b01000111100111011000: color_data = 12'b111011101110;
20'b01000111100111011001: color_data = 12'b111011101110;
20'b01000111100111011010: color_data = 12'b111011101110;
20'b01000111100111011011: color_data = 12'b111011101110;
20'b01000111100111011100: color_data = 12'b111011101110;
20'b01000111100111011110: color_data = 12'b111011101110;
20'b01000111100111011111: color_data = 12'b111011101110;
20'b01000111100111100000: color_data = 12'b111011101110;
20'b01000111100111100001: color_data = 12'b111011101110;
20'b01000111100111100010: color_data = 12'b111011101110;
20'b01000111100111100011: color_data = 12'b111011101110;
20'b01000111100111100100: color_data = 12'b111011101110;
20'b01000111100111100101: color_data = 12'b111011101110;
20'b01000111100111100110: color_data = 12'b111011101110;
20'b01000111100111100111: color_data = 12'b111011101110;
20'b01000111110010010110: color_data = 12'b111011101110;
20'b01000111110010010111: color_data = 12'b111011101110;
20'b01000111110010011000: color_data = 12'b111011101110;
20'b01000111110010011001: color_data = 12'b111011101110;
20'b01000111110010011010: color_data = 12'b111011101110;
20'b01000111110010011011: color_data = 12'b111011101110;
20'b01000111110010011100: color_data = 12'b111011101110;
20'b01000111110010011101: color_data = 12'b111011101110;
20'b01000111110010011110: color_data = 12'b111011101110;
20'b01000111110010011111: color_data = 12'b111011101110;
20'b01000111110010100001: color_data = 12'b111011101110;
20'b01000111110010100010: color_data = 12'b111011101110;
20'b01000111110010100011: color_data = 12'b111011101110;
20'b01000111110010100100: color_data = 12'b111011101110;
20'b01000111110010100101: color_data = 12'b111011101110;
20'b01000111110010100110: color_data = 12'b111011101110;
20'b01000111110010100111: color_data = 12'b111011101110;
20'b01000111110010101000: color_data = 12'b111011101110;
20'b01000111110010101001: color_data = 12'b111011101110;
20'b01000111110010101010: color_data = 12'b111011101110;
20'b01000111110011001101: color_data = 12'b111011101110;
20'b01000111110011001110: color_data = 12'b111011101110;
20'b01000111110011001111: color_data = 12'b111011101110;
20'b01000111110011010000: color_data = 12'b111011101110;
20'b01000111110011010001: color_data = 12'b111011101110;
20'b01000111110011010010: color_data = 12'b111011101110;
20'b01000111110011010011: color_data = 12'b111011101110;
20'b01000111110011010100: color_data = 12'b111011101110;
20'b01000111110011010101: color_data = 12'b111011101110;
20'b01000111110011010110: color_data = 12'b111011101110;
20'b01000111110011011000: color_data = 12'b111011101110;
20'b01000111110011011001: color_data = 12'b111011101110;
20'b01000111110011011010: color_data = 12'b111011101110;
20'b01000111110011011011: color_data = 12'b111011101110;
20'b01000111110011011100: color_data = 12'b111011101110;
20'b01000111110011011101: color_data = 12'b111011101110;
20'b01000111110011011110: color_data = 12'b111011101110;
20'b01000111110011011111: color_data = 12'b111011101110;
20'b01000111110011100000: color_data = 12'b111011101110;
20'b01000111110011100001: color_data = 12'b111011101110;
20'b01000111110011101101: color_data = 12'b111011101110;
20'b01000111110011101110: color_data = 12'b111011101110;
20'b01000111110011101111: color_data = 12'b111011101110;
20'b01000111110011110000: color_data = 12'b111011101110;
20'b01000111110011110001: color_data = 12'b111011101110;
20'b01000111110011110010: color_data = 12'b111011101110;
20'b01000111110011110011: color_data = 12'b111011101110;
20'b01000111110011110100: color_data = 12'b111011101110;
20'b01000111110011110101: color_data = 12'b111011101110;
20'b01000111110011110110: color_data = 12'b111011101110;
20'b01000111110011111000: color_data = 12'b111011101110;
20'b01000111110011111001: color_data = 12'b111011101110;
20'b01000111110011111010: color_data = 12'b111011101110;
20'b01000111110011111011: color_data = 12'b111011101110;
20'b01000111110011111100: color_data = 12'b111011101110;
20'b01000111110011111101: color_data = 12'b111011101110;
20'b01000111110011111110: color_data = 12'b111011101110;
20'b01000111110011111111: color_data = 12'b111011101110;
20'b01000111110100000000: color_data = 12'b111011101110;
20'b01000111110100000001: color_data = 12'b111011101110;
20'b01000111110100100100: color_data = 12'b111011101110;
20'b01000111110100100101: color_data = 12'b111011101110;
20'b01000111110100100110: color_data = 12'b111011101110;
20'b01000111110100100111: color_data = 12'b111011101110;
20'b01000111110100101000: color_data = 12'b111011101110;
20'b01000111110100101001: color_data = 12'b111011101110;
20'b01000111110100101010: color_data = 12'b111011101110;
20'b01000111110100101011: color_data = 12'b111011101110;
20'b01000111110100101100: color_data = 12'b111011101110;
20'b01000111110100101101: color_data = 12'b111011101110;
20'b01000111110100101111: color_data = 12'b111011101110;
20'b01000111110100110000: color_data = 12'b111011101110;
20'b01000111110100110001: color_data = 12'b111011101110;
20'b01000111110100110010: color_data = 12'b111011101110;
20'b01000111110100110011: color_data = 12'b111011101110;
20'b01000111110100110100: color_data = 12'b111011101110;
20'b01000111110100110101: color_data = 12'b111011101110;
20'b01000111110100110110: color_data = 12'b111011101110;
20'b01000111110100110111: color_data = 12'b111011101110;
20'b01000111110100111000: color_data = 12'b111011101110;
20'b01000111110101000100: color_data = 12'b111011101110;
20'b01000111110101000101: color_data = 12'b111011101110;
20'b01000111110101000110: color_data = 12'b111011101110;
20'b01000111110101000111: color_data = 12'b111011101110;
20'b01000111110101001000: color_data = 12'b111011101110;
20'b01000111110101001001: color_data = 12'b111011101110;
20'b01000111110101001010: color_data = 12'b111011101110;
20'b01000111110101001011: color_data = 12'b111011101110;
20'b01000111110101001100: color_data = 12'b111011101110;
20'b01000111110101001101: color_data = 12'b111011101110;
20'b01000111110101001111: color_data = 12'b111011101110;
20'b01000111110101010000: color_data = 12'b111011101110;
20'b01000111110101010001: color_data = 12'b111011101110;
20'b01000111110101010010: color_data = 12'b111011101110;
20'b01000111110101010011: color_data = 12'b111011101110;
20'b01000111110101010100: color_data = 12'b111011101110;
20'b01000111110101010101: color_data = 12'b111011101110;
20'b01000111110101010110: color_data = 12'b111011101110;
20'b01000111110101010111: color_data = 12'b111011101110;
20'b01000111110101011000: color_data = 12'b111011101110;
20'b01000111110110011100: color_data = 12'b111011101110;
20'b01000111110110011101: color_data = 12'b111011101110;
20'b01000111110110011110: color_data = 12'b111011101110;
20'b01000111110110011111: color_data = 12'b111011101110;
20'b01000111110110100000: color_data = 12'b111011101110;
20'b01000111110110100001: color_data = 12'b111011101110;
20'b01000111110110100010: color_data = 12'b111011101110;
20'b01000111110110100011: color_data = 12'b111011101110;
20'b01000111110110100100: color_data = 12'b111011101110;
20'b01000111110110100101: color_data = 12'b111011101110;
20'b01000111110110100111: color_data = 12'b111011101110;
20'b01000111110110101000: color_data = 12'b111011101110;
20'b01000111110110101001: color_data = 12'b111011101110;
20'b01000111110110101010: color_data = 12'b111011101110;
20'b01000111110110101011: color_data = 12'b111011101110;
20'b01000111110110101100: color_data = 12'b111011101110;
20'b01000111110110101101: color_data = 12'b111011101110;
20'b01000111110110101110: color_data = 12'b111011101110;
20'b01000111110110101111: color_data = 12'b111011101110;
20'b01000111110110110000: color_data = 12'b111011101110;
20'b01000111110111010011: color_data = 12'b111011101110;
20'b01000111110111010100: color_data = 12'b111011101110;
20'b01000111110111010101: color_data = 12'b111011101110;
20'b01000111110111010110: color_data = 12'b111011101110;
20'b01000111110111010111: color_data = 12'b111011101110;
20'b01000111110111011000: color_data = 12'b111011101110;
20'b01000111110111011001: color_data = 12'b111011101110;
20'b01000111110111011010: color_data = 12'b111011101110;
20'b01000111110111011011: color_data = 12'b111011101110;
20'b01000111110111011100: color_data = 12'b111011101110;
20'b01000111110111011110: color_data = 12'b111011101110;
20'b01000111110111011111: color_data = 12'b111011101110;
20'b01000111110111100000: color_data = 12'b111011101110;
20'b01000111110111100001: color_data = 12'b111011101110;
20'b01000111110111100010: color_data = 12'b111011101110;
20'b01000111110111100011: color_data = 12'b111011101110;
20'b01000111110111100100: color_data = 12'b111011101110;
20'b01000111110111100101: color_data = 12'b111011101110;
20'b01000111110111100110: color_data = 12'b111011101110;
20'b01000111110111100111: color_data = 12'b111011101110;
20'b01001000010010010110: color_data = 12'b111011101110;
20'b01001000010010010111: color_data = 12'b111011101110;
20'b01001000010010011000: color_data = 12'b111011101110;
20'b01001000010010011001: color_data = 12'b111011101110;
20'b01001000010010011010: color_data = 12'b111011101110;
20'b01001000010010011011: color_data = 12'b111011101110;
20'b01001000010010011100: color_data = 12'b111011101110;
20'b01001000010010011101: color_data = 12'b111011101110;
20'b01001000010010011110: color_data = 12'b111011101110;
20'b01001000010010011111: color_data = 12'b111011101110;
20'b01001000010010100001: color_data = 12'b111011101110;
20'b01001000010010100010: color_data = 12'b111011101110;
20'b01001000010010100011: color_data = 12'b111011101110;
20'b01001000010010100100: color_data = 12'b111011101110;
20'b01001000010010100101: color_data = 12'b111011101110;
20'b01001000010010100110: color_data = 12'b111011101110;
20'b01001000010010100111: color_data = 12'b111011101110;
20'b01001000010010101000: color_data = 12'b111011101110;
20'b01001000010010101001: color_data = 12'b111011101110;
20'b01001000010010101010: color_data = 12'b111011101110;
20'b01001000010011001101: color_data = 12'b111011101110;
20'b01001000010011001110: color_data = 12'b111011101110;
20'b01001000010011001111: color_data = 12'b111011101110;
20'b01001000010011010000: color_data = 12'b111011101110;
20'b01001000010011010001: color_data = 12'b111011101110;
20'b01001000010011010010: color_data = 12'b111011101110;
20'b01001000010011010011: color_data = 12'b111011101110;
20'b01001000010011010100: color_data = 12'b111011101110;
20'b01001000010011010101: color_data = 12'b111011101110;
20'b01001000010011010110: color_data = 12'b111011101110;
20'b01001000010011011000: color_data = 12'b111011101110;
20'b01001000010011011001: color_data = 12'b111011101110;
20'b01001000010011011010: color_data = 12'b111011101110;
20'b01001000010011011011: color_data = 12'b111011101110;
20'b01001000010011011100: color_data = 12'b111011101110;
20'b01001000010011011101: color_data = 12'b111011101110;
20'b01001000010011011110: color_data = 12'b111011101110;
20'b01001000010011011111: color_data = 12'b111011101110;
20'b01001000010011100000: color_data = 12'b111011101110;
20'b01001000010011100001: color_data = 12'b111011101110;
20'b01001000010011101101: color_data = 12'b111011101110;
20'b01001000010011101110: color_data = 12'b111011101110;
20'b01001000010011101111: color_data = 12'b111011101110;
20'b01001000010011110000: color_data = 12'b111011101110;
20'b01001000010011110001: color_data = 12'b111011101110;
20'b01001000010011110010: color_data = 12'b111011101110;
20'b01001000010011110011: color_data = 12'b111011101110;
20'b01001000010011110100: color_data = 12'b111011101110;
20'b01001000010011110101: color_data = 12'b111011101110;
20'b01001000010011110110: color_data = 12'b111011101110;
20'b01001000010011111000: color_data = 12'b111011101110;
20'b01001000010011111001: color_data = 12'b111011101110;
20'b01001000010011111010: color_data = 12'b111011101110;
20'b01001000010011111011: color_data = 12'b111011101110;
20'b01001000010011111100: color_data = 12'b111011101110;
20'b01001000010011111101: color_data = 12'b111011101110;
20'b01001000010011111110: color_data = 12'b111011101110;
20'b01001000010011111111: color_data = 12'b111011101110;
20'b01001000010100000000: color_data = 12'b111011101110;
20'b01001000010100000001: color_data = 12'b111011101110;
20'b01001000010100100100: color_data = 12'b111011101110;
20'b01001000010100100101: color_data = 12'b111011101110;
20'b01001000010100100110: color_data = 12'b111011101110;
20'b01001000010100100111: color_data = 12'b111011101110;
20'b01001000010100101000: color_data = 12'b111011101110;
20'b01001000010100101001: color_data = 12'b111011101110;
20'b01001000010100101010: color_data = 12'b111011101110;
20'b01001000010100101011: color_data = 12'b111011101110;
20'b01001000010100101100: color_data = 12'b111011101110;
20'b01001000010100101101: color_data = 12'b111011101110;
20'b01001000010100101111: color_data = 12'b111011101110;
20'b01001000010100110000: color_data = 12'b111011101110;
20'b01001000010100110001: color_data = 12'b111011101110;
20'b01001000010100110010: color_data = 12'b111011101110;
20'b01001000010100110011: color_data = 12'b111011101110;
20'b01001000010100110100: color_data = 12'b111011101110;
20'b01001000010100110101: color_data = 12'b111011101110;
20'b01001000010100110110: color_data = 12'b111011101110;
20'b01001000010100110111: color_data = 12'b111011101110;
20'b01001000010100111000: color_data = 12'b111011101110;
20'b01001000010101000100: color_data = 12'b111011101110;
20'b01001000010101000101: color_data = 12'b111011101110;
20'b01001000010101000110: color_data = 12'b111011101110;
20'b01001000010101000111: color_data = 12'b111011101110;
20'b01001000010101001000: color_data = 12'b111011101110;
20'b01001000010101001001: color_data = 12'b111011101110;
20'b01001000010101001010: color_data = 12'b111011101110;
20'b01001000010101001011: color_data = 12'b111011101110;
20'b01001000010101001100: color_data = 12'b111011101110;
20'b01001000010101001101: color_data = 12'b111011101110;
20'b01001000010101001111: color_data = 12'b111011101110;
20'b01001000010101010000: color_data = 12'b111011101110;
20'b01001000010101010001: color_data = 12'b111011101110;
20'b01001000010101010010: color_data = 12'b111011101110;
20'b01001000010101010011: color_data = 12'b111011101110;
20'b01001000010101010100: color_data = 12'b111011101110;
20'b01001000010101010101: color_data = 12'b111011101110;
20'b01001000010101010110: color_data = 12'b111011101110;
20'b01001000010101010111: color_data = 12'b111011101110;
20'b01001000010101011000: color_data = 12'b111011101110;
20'b01001000010101011010: color_data = 12'b111011101110;
20'b01001000010101011011: color_data = 12'b111011101110;
20'b01001000010101011100: color_data = 12'b111011101110;
20'b01001000010101011101: color_data = 12'b111011101110;
20'b01001000010101011110: color_data = 12'b111011101110;
20'b01001000010101011111: color_data = 12'b111011101110;
20'b01001000010101100000: color_data = 12'b111011101110;
20'b01001000010101100001: color_data = 12'b111011101110;
20'b01001000010101100010: color_data = 12'b111011101110;
20'b01001000010101100011: color_data = 12'b111011101110;
20'b01001000010101100101: color_data = 12'b111011101110;
20'b01001000010101100110: color_data = 12'b111011101110;
20'b01001000010101100111: color_data = 12'b111011101110;
20'b01001000010101101000: color_data = 12'b111011101110;
20'b01001000010101101001: color_data = 12'b111011101110;
20'b01001000010101101010: color_data = 12'b111011101110;
20'b01001000010101101011: color_data = 12'b111011101110;
20'b01001000010101101100: color_data = 12'b111011101110;
20'b01001000010101101101: color_data = 12'b111011101110;
20'b01001000010101101110: color_data = 12'b111011101110;
20'b01001000010101110000: color_data = 12'b111011101110;
20'b01001000010101110001: color_data = 12'b111011101110;
20'b01001000010101110010: color_data = 12'b111011101110;
20'b01001000010101110011: color_data = 12'b111011101110;
20'b01001000010101110100: color_data = 12'b111011101110;
20'b01001000010101110101: color_data = 12'b111011101110;
20'b01001000010101110110: color_data = 12'b111011101110;
20'b01001000010101110111: color_data = 12'b111011101110;
20'b01001000010101111000: color_data = 12'b111011101110;
20'b01001000010101111001: color_data = 12'b111011101110;
20'b01001000010110011100: color_data = 12'b111011101110;
20'b01001000010110011101: color_data = 12'b111011101110;
20'b01001000010110011110: color_data = 12'b111011101110;
20'b01001000010110011111: color_data = 12'b111011101110;
20'b01001000010110100000: color_data = 12'b111011101110;
20'b01001000010110100001: color_data = 12'b111011101110;
20'b01001000010110100010: color_data = 12'b111011101110;
20'b01001000010110100011: color_data = 12'b111011101110;
20'b01001000010110100100: color_data = 12'b111011101110;
20'b01001000010110100101: color_data = 12'b111011101110;
20'b01001000010110100111: color_data = 12'b111011101110;
20'b01001000010110101000: color_data = 12'b111011101110;
20'b01001000010110101001: color_data = 12'b111011101110;
20'b01001000010110101010: color_data = 12'b111011101110;
20'b01001000010110101011: color_data = 12'b111011101110;
20'b01001000010110101100: color_data = 12'b111011101110;
20'b01001000010110101101: color_data = 12'b111011101110;
20'b01001000010110101110: color_data = 12'b111011101110;
20'b01001000010110101111: color_data = 12'b111011101110;
20'b01001000010110110000: color_data = 12'b111011101110;
20'b01001000010110111101: color_data = 12'b111011101110;
20'b01001000010110111110: color_data = 12'b111011101110;
20'b01001000010110111111: color_data = 12'b111011101110;
20'b01001000010111000000: color_data = 12'b111011101110;
20'b01001000010111000001: color_data = 12'b111011101110;
20'b01001000010111000010: color_data = 12'b111011101110;
20'b01001000010111000011: color_data = 12'b111011101110;
20'b01001000010111000100: color_data = 12'b111011101110;
20'b01001000010111000101: color_data = 12'b111011101110;
20'b01001000010111000110: color_data = 12'b111011101110;
20'b01001000010111001000: color_data = 12'b111011101110;
20'b01001000010111001001: color_data = 12'b111011101110;
20'b01001000010111001010: color_data = 12'b111011101110;
20'b01001000010111001011: color_data = 12'b111011101110;
20'b01001000010111001100: color_data = 12'b111011101110;
20'b01001000010111001101: color_data = 12'b111011101110;
20'b01001000010111001110: color_data = 12'b111011101110;
20'b01001000010111001111: color_data = 12'b111011101110;
20'b01001000010111010000: color_data = 12'b111011101110;
20'b01001000010111010001: color_data = 12'b111011101110;
20'b01001000010111010011: color_data = 12'b111011101110;
20'b01001000010111010100: color_data = 12'b111011101110;
20'b01001000010111010101: color_data = 12'b111011101110;
20'b01001000010111010110: color_data = 12'b111011101110;
20'b01001000010111010111: color_data = 12'b111011101110;
20'b01001000010111011000: color_data = 12'b111011101110;
20'b01001000010111011001: color_data = 12'b111011101110;
20'b01001000010111011010: color_data = 12'b111011101110;
20'b01001000010111011011: color_data = 12'b111011101110;
20'b01001000010111011100: color_data = 12'b111011101110;
20'b01001000100010010110: color_data = 12'b111011101110;
20'b01001000100010010111: color_data = 12'b111011101110;
20'b01001000100010011000: color_data = 12'b111011101110;
20'b01001000100010011001: color_data = 12'b111011101110;
20'b01001000100010011010: color_data = 12'b111011101110;
20'b01001000100010011011: color_data = 12'b111011101110;
20'b01001000100010011100: color_data = 12'b111011101110;
20'b01001000100010011101: color_data = 12'b111011101110;
20'b01001000100010011110: color_data = 12'b111011101110;
20'b01001000100010011111: color_data = 12'b111011101110;
20'b01001000100010100001: color_data = 12'b111011101110;
20'b01001000100010100010: color_data = 12'b111011101110;
20'b01001000100010100011: color_data = 12'b111011101110;
20'b01001000100010100100: color_data = 12'b111011101110;
20'b01001000100010100101: color_data = 12'b111011101110;
20'b01001000100010100110: color_data = 12'b111011101110;
20'b01001000100010100111: color_data = 12'b111011101110;
20'b01001000100010101000: color_data = 12'b111011101110;
20'b01001000100010101001: color_data = 12'b111011101110;
20'b01001000100010101010: color_data = 12'b111011101110;
20'b01001000100011001101: color_data = 12'b111011101110;
20'b01001000100011001110: color_data = 12'b111011101110;
20'b01001000100011001111: color_data = 12'b111011101110;
20'b01001000100011010000: color_data = 12'b111011101110;
20'b01001000100011010001: color_data = 12'b111011101110;
20'b01001000100011010010: color_data = 12'b111011101110;
20'b01001000100011010011: color_data = 12'b111011101110;
20'b01001000100011010100: color_data = 12'b111011101110;
20'b01001000100011010101: color_data = 12'b111011101110;
20'b01001000100011010110: color_data = 12'b111011101110;
20'b01001000100011011000: color_data = 12'b111011101110;
20'b01001000100011011001: color_data = 12'b111011101110;
20'b01001000100011011010: color_data = 12'b111011101110;
20'b01001000100011011011: color_data = 12'b111011101110;
20'b01001000100011011100: color_data = 12'b111011101110;
20'b01001000100011011101: color_data = 12'b111011101110;
20'b01001000100011011110: color_data = 12'b111011101110;
20'b01001000100011011111: color_data = 12'b111011101110;
20'b01001000100011100000: color_data = 12'b111011101110;
20'b01001000100011100001: color_data = 12'b111011101110;
20'b01001000100011101101: color_data = 12'b111011101110;
20'b01001000100011101110: color_data = 12'b111011101110;
20'b01001000100011101111: color_data = 12'b111011101110;
20'b01001000100011110000: color_data = 12'b111011101110;
20'b01001000100011110001: color_data = 12'b111011101110;
20'b01001000100011110010: color_data = 12'b111011101110;
20'b01001000100011110011: color_data = 12'b111011101110;
20'b01001000100011110100: color_data = 12'b111011101110;
20'b01001000100011110101: color_data = 12'b111011101110;
20'b01001000100011110110: color_data = 12'b111011101110;
20'b01001000100011111000: color_data = 12'b111011101110;
20'b01001000100011111001: color_data = 12'b111011101110;
20'b01001000100011111010: color_data = 12'b111011101110;
20'b01001000100011111011: color_data = 12'b111011101110;
20'b01001000100011111100: color_data = 12'b111011101110;
20'b01001000100011111101: color_data = 12'b111011101110;
20'b01001000100011111110: color_data = 12'b111011101110;
20'b01001000100011111111: color_data = 12'b111011101110;
20'b01001000100100000000: color_data = 12'b111011101110;
20'b01001000100100000001: color_data = 12'b111011101110;
20'b01001000100100100100: color_data = 12'b111011101110;
20'b01001000100100100101: color_data = 12'b111011101110;
20'b01001000100100100110: color_data = 12'b111011101110;
20'b01001000100100100111: color_data = 12'b111011101110;
20'b01001000100100101000: color_data = 12'b111011101110;
20'b01001000100100101001: color_data = 12'b111011101110;
20'b01001000100100101010: color_data = 12'b111011101110;
20'b01001000100100101011: color_data = 12'b111011101110;
20'b01001000100100101100: color_data = 12'b111011101110;
20'b01001000100100101101: color_data = 12'b111011101110;
20'b01001000100100101111: color_data = 12'b111011101110;
20'b01001000100100110000: color_data = 12'b111011101110;
20'b01001000100100110001: color_data = 12'b111011101110;
20'b01001000100100110010: color_data = 12'b111011101110;
20'b01001000100100110011: color_data = 12'b111011101110;
20'b01001000100100110100: color_data = 12'b111011101110;
20'b01001000100100110101: color_data = 12'b111011101110;
20'b01001000100100110110: color_data = 12'b111011101110;
20'b01001000100100110111: color_data = 12'b111011101110;
20'b01001000100100111000: color_data = 12'b111011101110;
20'b01001000100101000100: color_data = 12'b111011101110;
20'b01001000100101000101: color_data = 12'b111011101110;
20'b01001000100101000110: color_data = 12'b111011101110;
20'b01001000100101000111: color_data = 12'b111011101110;
20'b01001000100101001000: color_data = 12'b111011101110;
20'b01001000100101001001: color_data = 12'b111011101110;
20'b01001000100101001010: color_data = 12'b111011101110;
20'b01001000100101001011: color_data = 12'b111011101110;
20'b01001000100101001100: color_data = 12'b111011101110;
20'b01001000100101001101: color_data = 12'b111011101110;
20'b01001000100101001111: color_data = 12'b111011101110;
20'b01001000100101010000: color_data = 12'b111011101110;
20'b01001000100101010001: color_data = 12'b111011101110;
20'b01001000100101010010: color_data = 12'b111011101110;
20'b01001000100101010011: color_data = 12'b111011101110;
20'b01001000100101010100: color_data = 12'b111011101110;
20'b01001000100101010101: color_data = 12'b111011101110;
20'b01001000100101010110: color_data = 12'b111011101110;
20'b01001000100101010111: color_data = 12'b111011101110;
20'b01001000100101011000: color_data = 12'b111011101110;
20'b01001000100101011010: color_data = 12'b111011101110;
20'b01001000100101011011: color_data = 12'b111011101110;
20'b01001000100101011100: color_data = 12'b111011101110;
20'b01001000100101011101: color_data = 12'b111011101110;
20'b01001000100101011110: color_data = 12'b111011101110;
20'b01001000100101011111: color_data = 12'b111011101110;
20'b01001000100101100000: color_data = 12'b111011101110;
20'b01001000100101100001: color_data = 12'b111011101110;
20'b01001000100101100010: color_data = 12'b111011101110;
20'b01001000100101100011: color_data = 12'b111011101110;
20'b01001000100101100101: color_data = 12'b111011101110;
20'b01001000100101100110: color_data = 12'b111011101110;
20'b01001000100101100111: color_data = 12'b111011101110;
20'b01001000100101101000: color_data = 12'b111011101110;
20'b01001000100101101001: color_data = 12'b111011101110;
20'b01001000100101101010: color_data = 12'b111011101110;
20'b01001000100101101011: color_data = 12'b111011101110;
20'b01001000100101101100: color_data = 12'b111011101110;
20'b01001000100101101101: color_data = 12'b111011101110;
20'b01001000100101101110: color_data = 12'b111011101110;
20'b01001000100101110000: color_data = 12'b111011101110;
20'b01001000100101110001: color_data = 12'b111011101110;
20'b01001000100101110010: color_data = 12'b111011101110;
20'b01001000100101110011: color_data = 12'b111011101110;
20'b01001000100101110100: color_data = 12'b111011101110;
20'b01001000100101110101: color_data = 12'b111011101110;
20'b01001000100101110110: color_data = 12'b111011101110;
20'b01001000100101110111: color_data = 12'b111011101110;
20'b01001000100101111000: color_data = 12'b111011101110;
20'b01001000100101111001: color_data = 12'b111011101110;
20'b01001000100110011100: color_data = 12'b111011101110;
20'b01001000100110011101: color_data = 12'b111011101110;
20'b01001000100110011110: color_data = 12'b111011101110;
20'b01001000100110011111: color_data = 12'b111011101110;
20'b01001000100110100000: color_data = 12'b111011101110;
20'b01001000100110100001: color_data = 12'b111011101110;
20'b01001000100110100010: color_data = 12'b111011101110;
20'b01001000100110100011: color_data = 12'b111011101110;
20'b01001000100110100100: color_data = 12'b111011101110;
20'b01001000100110100101: color_data = 12'b111011101110;
20'b01001000100110100111: color_data = 12'b111011101110;
20'b01001000100110101000: color_data = 12'b111011101110;
20'b01001000100110101001: color_data = 12'b111011101110;
20'b01001000100110101010: color_data = 12'b111011101110;
20'b01001000100110101011: color_data = 12'b111011101110;
20'b01001000100110101100: color_data = 12'b111011101110;
20'b01001000100110101101: color_data = 12'b111011101110;
20'b01001000100110101110: color_data = 12'b111011101110;
20'b01001000100110101111: color_data = 12'b111011101110;
20'b01001000100110110000: color_data = 12'b111011101110;
20'b01001000100110111101: color_data = 12'b111011101110;
20'b01001000100110111110: color_data = 12'b111011101110;
20'b01001000100110111111: color_data = 12'b111011101110;
20'b01001000100111000000: color_data = 12'b111011101110;
20'b01001000100111000001: color_data = 12'b111011101110;
20'b01001000100111000010: color_data = 12'b111011101110;
20'b01001000100111000011: color_data = 12'b111011101110;
20'b01001000100111000100: color_data = 12'b111011101110;
20'b01001000100111000101: color_data = 12'b111011101110;
20'b01001000100111000110: color_data = 12'b111011101110;
20'b01001000100111001000: color_data = 12'b111011101110;
20'b01001000100111001001: color_data = 12'b111011101110;
20'b01001000100111001010: color_data = 12'b111011101110;
20'b01001000100111001011: color_data = 12'b111011101110;
20'b01001000100111001100: color_data = 12'b111011101110;
20'b01001000100111001101: color_data = 12'b111011101110;
20'b01001000100111001110: color_data = 12'b111011101110;
20'b01001000100111001111: color_data = 12'b111011101110;
20'b01001000100111010000: color_data = 12'b111011101110;
20'b01001000100111010001: color_data = 12'b111011101110;
20'b01001000100111010011: color_data = 12'b111011101110;
20'b01001000100111010100: color_data = 12'b111011101110;
20'b01001000100111010101: color_data = 12'b111011101110;
20'b01001000100111010110: color_data = 12'b111011101110;
20'b01001000100111010111: color_data = 12'b111011101110;
20'b01001000100111011000: color_data = 12'b111011101110;
20'b01001000100111011001: color_data = 12'b111011101110;
20'b01001000100111011010: color_data = 12'b111011101110;
20'b01001000100111011011: color_data = 12'b111011101110;
20'b01001000100111011100: color_data = 12'b111011101110;
20'b01001000110010010110: color_data = 12'b111011101110;
20'b01001000110010010111: color_data = 12'b111011101110;
20'b01001000110010011000: color_data = 12'b111011101110;
20'b01001000110010011001: color_data = 12'b111011101110;
20'b01001000110010011010: color_data = 12'b111011101110;
20'b01001000110010011011: color_data = 12'b111011101110;
20'b01001000110010011100: color_data = 12'b111011101110;
20'b01001000110010011101: color_data = 12'b111011101110;
20'b01001000110010011110: color_data = 12'b111011101110;
20'b01001000110010011111: color_data = 12'b111011101110;
20'b01001000110010100001: color_data = 12'b111011101110;
20'b01001000110010100010: color_data = 12'b111011101110;
20'b01001000110010100011: color_data = 12'b111011101110;
20'b01001000110010100100: color_data = 12'b111011101110;
20'b01001000110010100101: color_data = 12'b111011101110;
20'b01001000110010100110: color_data = 12'b111011101110;
20'b01001000110010100111: color_data = 12'b111011101110;
20'b01001000110010101000: color_data = 12'b111011101110;
20'b01001000110010101001: color_data = 12'b111011101110;
20'b01001000110010101010: color_data = 12'b111011101110;
20'b01001000110011001101: color_data = 12'b111011101110;
20'b01001000110011001110: color_data = 12'b111011101110;
20'b01001000110011001111: color_data = 12'b111011101110;
20'b01001000110011010000: color_data = 12'b111011101110;
20'b01001000110011010001: color_data = 12'b111011101110;
20'b01001000110011010010: color_data = 12'b111011101110;
20'b01001000110011010011: color_data = 12'b111011101110;
20'b01001000110011010100: color_data = 12'b111011101110;
20'b01001000110011010101: color_data = 12'b111011101110;
20'b01001000110011010110: color_data = 12'b111011101110;
20'b01001000110011011000: color_data = 12'b111011101110;
20'b01001000110011011001: color_data = 12'b111011101110;
20'b01001000110011011010: color_data = 12'b111011101110;
20'b01001000110011011011: color_data = 12'b111011101110;
20'b01001000110011011100: color_data = 12'b111011101110;
20'b01001000110011011101: color_data = 12'b111011101110;
20'b01001000110011011110: color_data = 12'b111011101110;
20'b01001000110011011111: color_data = 12'b111011101110;
20'b01001000110011100000: color_data = 12'b111011101110;
20'b01001000110011100001: color_data = 12'b111011101110;
20'b01001000110011101101: color_data = 12'b111011101110;
20'b01001000110011101110: color_data = 12'b111011101110;
20'b01001000110011101111: color_data = 12'b111011101110;
20'b01001000110011110000: color_data = 12'b111011101110;
20'b01001000110011110001: color_data = 12'b111011101110;
20'b01001000110011110010: color_data = 12'b111011101110;
20'b01001000110011110011: color_data = 12'b111011101110;
20'b01001000110011110100: color_data = 12'b111011101110;
20'b01001000110011110101: color_data = 12'b111011101110;
20'b01001000110011110110: color_data = 12'b111011101110;
20'b01001000110011111000: color_data = 12'b111011101110;
20'b01001000110011111001: color_data = 12'b111011101110;
20'b01001000110011111010: color_data = 12'b111011101110;
20'b01001000110011111011: color_data = 12'b111011101110;
20'b01001000110011111100: color_data = 12'b111011101110;
20'b01001000110011111101: color_data = 12'b111011101110;
20'b01001000110011111110: color_data = 12'b111011101110;
20'b01001000110011111111: color_data = 12'b111011101110;
20'b01001000110100000000: color_data = 12'b111011101110;
20'b01001000110100000001: color_data = 12'b111011101110;
20'b01001000110100100100: color_data = 12'b111011101110;
20'b01001000110100100101: color_data = 12'b111011101110;
20'b01001000110100100110: color_data = 12'b111011101110;
20'b01001000110100100111: color_data = 12'b111011101110;
20'b01001000110100101000: color_data = 12'b111011101110;
20'b01001000110100101001: color_data = 12'b111011101110;
20'b01001000110100101010: color_data = 12'b111011101110;
20'b01001000110100101011: color_data = 12'b111011101110;
20'b01001000110100101100: color_data = 12'b111011101110;
20'b01001000110100101101: color_data = 12'b111011101110;
20'b01001000110100101111: color_data = 12'b111011101110;
20'b01001000110100110000: color_data = 12'b111011101110;
20'b01001000110100110001: color_data = 12'b111011101110;
20'b01001000110100110010: color_data = 12'b111011101110;
20'b01001000110100110011: color_data = 12'b111011101110;
20'b01001000110100110100: color_data = 12'b111011101110;
20'b01001000110100110101: color_data = 12'b111011101110;
20'b01001000110100110110: color_data = 12'b111011101110;
20'b01001000110100110111: color_data = 12'b111011101110;
20'b01001000110100111000: color_data = 12'b111011101110;
20'b01001000110101000100: color_data = 12'b111011101110;
20'b01001000110101000101: color_data = 12'b111011101110;
20'b01001000110101000110: color_data = 12'b111011101110;
20'b01001000110101000111: color_data = 12'b111011101110;
20'b01001000110101001000: color_data = 12'b111011101110;
20'b01001000110101001001: color_data = 12'b111011101110;
20'b01001000110101001010: color_data = 12'b111011101110;
20'b01001000110101001011: color_data = 12'b111011101110;
20'b01001000110101001100: color_data = 12'b111011101110;
20'b01001000110101001101: color_data = 12'b111011101110;
20'b01001000110101001111: color_data = 12'b111011101110;
20'b01001000110101010000: color_data = 12'b111011101110;
20'b01001000110101010001: color_data = 12'b111011101110;
20'b01001000110101010010: color_data = 12'b111011101110;
20'b01001000110101010011: color_data = 12'b111011101110;
20'b01001000110101010100: color_data = 12'b111011101110;
20'b01001000110101010101: color_data = 12'b111011101110;
20'b01001000110101010110: color_data = 12'b111011101110;
20'b01001000110101010111: color_data = 12'b111011101110;
20'b01001000110101011000: color_data = 12'b111011101110;
20'b01001000110101011010: color_data = 12'b111011101110;
20'b01001000110101011011: color_data = 12'b111011101110;
20'b01001000110101011100: color_data = 12'b111011101110;
20'b01001000110101011101: color_data = 12'b111011101110;
20'b01001000110101011110: color_data = 12'b111011101110;
20'b01001000110101011111: color_data = 12'b111011101110;
20'b01001000110101100000: color_data = 12'b111011101110;
20'b01001000110101100001: color_data = 12'b111011101110;
20'b01001000110101100010: color_data = 12'b111011101110;
20'b01001000110101100011: color_data = 12'b111011101110;
20'b01001000110101100101: color_data = 12'b111011101110;
20'b01001000110101100110: color_data = 12'b111011101110;
20'b01001000110101100111: color_data = 12'b111011101110;
20'b01001000110101101000: color_data = 12'b111011101110;
20'b01001000110101101001: color_data = 12'b111011101110;
20'b01001000110101101010: color_data = 12'b111011101110;
20'b01001000110101101011: color_data = 12'b111011101110;
20'b01001000110101101100: color_data = 12'b111011101110;
20'b01001000110101101101: color_data = 12'b111011101110;
20'b01001000110101101110: color_data = 12'b111011101110;
20'b01001000110101110000: color_data = 12'b111011101110;
20'b01001000110101110001: color_data = 12'b111011101110;
20'b01001000110101110010: color_data = 12'b111011101110;
20'b01001000110101110011: color_data = 12'b111011101110;
20'b01001000110101110100: color_data = 12'b111011101110;
20'b01001000110101110101: color_data = 12'b111011101110;
20'b01001000110101110110: color_data = 12'b111011101110;
20'b01001000110101110111: color_data = 12'b111011101110;
20'b01001000110101111000: color_data = 12'b111011101110;
20'b01001000110101111001: color_data = 12'b111011101110;
20'b01001000110110011100: color_data = 12'b111011101110;
20'b01001000110110011101: color_data = 12'b111011101110;
20'b01001000110110011110: color_data = 12'b111011101110;
20'b01001000110110011111: color_data = 12'b111011101110;
20'b01001000110110100000: color_data = 12'b111011101110;
20'b01001000110110100001: color_data = 12'b111011101110;
20'b01001000110110100010: color_data = 12'b111011101110;
20'b01001000110110100011: color_data = 12'b111011101110;
20'b01001000110110100100: color_data = 12'b111011101110;
20'b01001000110110100101: color_data = 12'b111011101110;
20'b01001000110110100111: color_data = 12'b111011101110;
20'b01001000110110101000: color_data = 12'b111011101110;
20'b01001000110110101001: color_data = 12'b111011101110;
20'b01001000110110101010: color_data = 12'b111011101110;
20'b01001000110110101011: color_data = 12'b111011101110;
20'b01001000110110101100: color_data = 12'b111011101110;
20'b01001000110110101101: color_data = 12'b111011101110;
20'b01001000110110101110: color_data = 12'b111011101110;
20'b01001000110110101111: color_data = 12'b111011101110;
20'b01001000110110110000: color_data = 12'b111011101110;
20'b01001000110110111101: color_data = 12'b111011101110;
20'b01001000110110111110: color_data = 12'b111011101110;
20'b01001000110110111111: color_data = 12'b111011101110;
20'b01001000110111000000: color_data = 12'b111011101110;
20'b01001000110111000001: color_data = 12'b111011101110;
20'b01001000110111000010: color_data = 12'b111011101110;
20'b01001000110111000011: color_data = 12'b111011101110;
20'b01001000110111000100: color_data = 12'b111011101110;
20'b01001000110111000101: color_data = 12'b111011101110;
20'b01001000110111000110: color_data = 12'b111011101110;
20'b01001000110111001000: color_data = 12'b111011101110;
20'b01001000110111001001: color_data = 12'b111011101110;
20'b01001000110111001010: color_data = 12'b111011101110;
20'b01001000110111001011: color_data = 12'b111011101110;
20'b01001000110111001100: color_data = 12'b111011101110;
20'b01001000110111001101: color_data = 12'b111011101110;
20'b01001000110111001110: color_data = 12'b111011101110;
20'b01001000110111001111: color_data = 12'b111011101110;
20'b01001000110111010000: color_data = 12'b111011101110;
20'b01001000110111010001: color_data = 12'b111011101110;
20'b01001000110111010011: color_data = 12'b111011101110;
20'b01001000110111010100: color_data = 12'b111011101110;
20'b01001000110111010101: color_data = 12'b111011101110;
20'b01001000110111010110: color_data = 12'b111011101110;
20'b01001000110111010111: color_data = 12'b111011101110;
20'b01001000110111011000: color_data = 12'b111011101110;
20'b01001000110111011001: color_data = 12'b111011101110;
20'b01001000110111011010: color_data = 12'b111011101110;
20'b01001000110111011011: color_data = 12'b111011101110;
20'b01001000110111011100: color_data = 12'b111011101110;
20'b01001001000010010110: color_data = 12'b111011101110;
20'b01001001000010010111: color_data = 12'b111011101110;
20'b01001001000010011000: color_data = 12'b111011101110;
20'b01001001000010011001: color_data = 12'b111011101110;
20'b01001001000010011010: color_data = 12'b111011101110;
20'b01001001000010011011: color_data = 12'b111011101110;
20'b01001001000010011100: color_data = 12'b111011101110;
20'b01001001000010011101: color_data = 12'b111011101110;
20'b01001001000010011110: color_data = 12'b111011101110;
20'b01001001000010011111: color_data = 12'b111011101110;
20'b01001001000010100001: color_data = 12'b111011101110;
20'b01001001000010100010: color_data = 12'b111011101110;
20'b01001001000010100011: color_data = 12'b111011101110;
20'b01001001000010100100: color_data = 12'b111011101110;
20'b01001001000010100101: color_data = 12'b111011101110;
20'b01001001000010100110: color_data = 12'b111011101110;
20'b01001001000010100111: color_data = 12'b111011101110;
20'b01001001000010101000: color_data = 12'b111011101110;
20'b01001001000010101001: color_data = 12'b111011101110;
20'b01001001000010101010: color_data = 12'b111011101110;
20'b01001001000011001101: color_data = 12'b111011101110;
20'b01001001000011001110: color_data = 12'b111011101110;
20'b01001001000011001111: color_data = 12'b111011101110;
20'b01001001000011010000: color_data = 12'b111011101110;
20'b01001001000011010001: color_data = 12'b111011101110;
20'b01001001000011010010: color_data = 12'b111011101110;
20'b01001001000011010011: color_data = 12'b111011101110;
20'b01001001000011010100: color_data = 12'b111011101110;
20'b01001001000011010101: color_data = 12'b111011101110;
20'b01001001000011010110: color_data = 12'b111011101110;
20'b01001001000011011000: color_data = 12'b111011101110;
20'b01001001000011011001: color_data = 12'b111011101110;
20'b01001001000011011010: color_data = 12'b111011101110;
20'b01001001000011011011: color_data = 12'b111011101110;
20'b01001001000011011100: color_data = 12'b111011101110;
20'b01001001000011011101: color_data = 12'b111011101110;
20'b01001001000011011110: color_data = 12'b111011101110;
20'b01001001000011011111: color_data = 12'b111011101110;
20'b01001001000011100000: color_data = 12'b111011101110;
20'b01001001000011100001: color_data = 12'b111011101110;
20'b01001001000011101101: color_data = 12'b111011101110;
20'b01001001000011101110: color_data = 12'b111011101110;
20'b01001001000011101111: color_data = 12'b111011101110;
20'b01001001000011110000: color_data = 12'b111011101110;
20'b01001001000011110001: color_data = 12'b111011101110;
20'b01001001000011110010: color_data = 12'b111011101110;
20'b01001001000011110011: color_data = 12'b111011101110;
20'b01001001000011110100: color_data = 12'b111011101110;
20'b01001001000011110101: color_data = 12'b111011101110;
20'b01001001000011110110: color_data = 12'b111011101110;
20'b01001001000011111000: color_data = 12'b111011101110;
20'b01001001000011111001: color_data = 12'b111011101110;
20'b01001001000011111010: color_data = 12'b111011101110;
20'b01001001000011111011: color_data = 12'b111011101110;
20'b01001001000011111100: color_data = 12'b111011101110;
20'b01001001000011111101: color_data = 12'b111011101110;
20'b01001001000011111110: color_data = 12'b111011101110;
20'b01001001000011111111: color_data = 12'b111011101110;
20'b01001001000100000000: color_data = 12'b111011101110;
20'b01001001000100000001: color_data = 12'b111011101110;
20'b01001001000100100100: color_data = 12'b111011101110;
20'b01001001000100100101: color_data = 12'b111011101110;
20'b01001001000100100110: color_data = 12'b111011101110;
20'b01001001000100100111: color_data = 12'b111011101110;
20'b01001001000100101000: color_data = 12'b111011101110;
20'b01001001000100101001: color_data = 12'b111011101110;
20'b01001001000100101010: color_data = 12'b111011101110;
20'b01001001000100101011: color_data = 12'b111011101110;
20'b01001001000100101100: color_data = 12'b111011101110;
20'b01001001000100101101: color_data = 12'b111011101110;
20'b01001001000100101111: color_data = 12'b111011101110;
20'b01001001000100110000: color_data = 12'b111011101110;
20'b01001001000100110001: color_data = 12'b111011101110;
20'b01001001000100110010: color_data = 12'b111011101110;
20'b01001001000100110011: color_data = 12'b111011101110;
20'b01001001000100110100: color_data = 12'b111011101110;
20'b01001001000100110101: color_data = 12'b111011101110;
20'b01001001000100110110: color_data = 12'b111011101110;
20'b01001001000100110111: color_data = 12'b111011101110;
20'b01001001000100111000: color_data = 12'b111011101110;
20'b01001001000101000100: color_data = 12'b111011101110;
20'b01001001000101000101: color_data = 12'b111011101110;
20'b01001001000101000110: color_data = 12'b111011101110;
20'b01001001000101000111: color_data = 12'b111011101110;
20'b01001001000101001000: color_data = 12'b111011101110;
20'b01001001000101001001: color_data = 12'b111011101110;
20'b01001001000101001010: color_data = 12'b111011101110;
20'b01001001000101001011: color_data = 12'b111011101110;
20'b01001001000101001100: color_data = 12'b111011101110;
20'b01001001000101001101: color_data = 12'b111011101110;
20'b01001001000101001111: color_data = 12'b111011101110;
20'b01001001000101010000: color_data = 12'b111011101110;
20'b01001001000101010001: color_data = 12'b111011101110;
20'b01001001000101010010: color_data = 12'b111011101110;
20'b01001001000101010011: color_data = 12'b111011101110;
20'b01001001000101010100: color_data = 12'b111011101110;
20'b01001001000101010101: color_data = 12'b111011101110;
20'b01001001000101010110: color_data = 12'b111011101110;
20'b01001001000101010111: color_data = 12'b111011101110;
20'b01001001000101011000: color_data = 12'b111011101110;
20'b01001001000101011010: color_data = 12'b111011101110;
20'b01001001000101011011: color_data = 12'b111011101110;
20'b01001001000101011100: color_data = 12'b111011101110;
20'b01001001000101011101: color_data = 12'b111011101110;
20'b01001001000101011110: color_data = 12'b111011101110;
20'b01001001000101011111: color_data = 12'b111011101110;
20'b01001001000101100000: color_data = 12'b111011101110;
20'b01001001000101100001: color_data = 12'b111011101110;
20'b01001001000101100010: color_data = 12'b111011101110;
20'b01001001000101100011: color_data = 12'b111011101110;
20'b01001001000101100101: color_data = 12'b111011101110;
20'b01001001000101100110: color_data = 12'b111011101110;
20'b01001001000101100111: color_data = 12'b111011101110;
20'b01001001000101101000: color_data = 12'b111011101110;
20'b01001001000101101001: color_data = 12'b111011101110;
20'b01001001000101101010: color_data = 12'b111011101110;
20'b01001001000101101011: color_data = 12'b111011101110;
20'b01001001000101101100: color_data = 12'b111011101110;
20'b01001001000101101101: color_data = 12'b111011101110;
20'b01001001000101101110: color_data = 12'b111011101110;
20'b01001001000101110000: color_data = 12'b111011101110;
20'b01001001000101110001: color_data = 12'b111011101110;
20'b01001001000101110010: color_data = 12'b111011101110;
20'b01001001000101110011: color_data = 12'b111011101110;
20'b01001001000101110100: color_data = 12'b111011101110;
20'b01001001000101110101: color_data = 12'b111011101110;
20'b01001001000101110110: color_data = 12'b111011101110;
20'b01001001000101110111: color_data = 12'b111011101110;
20'b01001001000101111000: color_data = 12'b111011101110;
20'b01001001000101111001: color_data = 12'b111011101110;
20'b01001001000110011100: color_data = 12'b111011101110;
20'b01001001000110011101: color_data = 12'b111011101110;
20'b01001001000110011110: color_data = 12'b111011101110;
20'b01001001000110011111: color_data = 12'b111011101110;
20'b01001001000110100000: color_data = 12'b111011101110;
20'b01001001000110100001: color_data = 12'b111011101110;
20'b01001001000110100010: color_data = 12'b111011101110;
20'b01001001000110100011: color_data = 12'b111011101110;
20'b01001001000110100100: color_data = 12'b111011101110;
20'b01001001000110100101: color_data = 12'b111011101110;
20'b01001001000110100111: color_data = 12'b111011101110;
20'b01001001000110101000: color_data = 12'b111011101110;
20'b01001001000110101001: color_data = 12'b111011101110;
20'b01001001000110101010: color_data = 12'b111011101110;
20'b01001001000110101011: color_data = 12'b111011101110;
20'b01001001000110101100: color_data = 12'b111011101110;
20'b01001001000110101101: color_data = 12'b111011101110;
20'b01001001000110101110: color_data = 12'b111011101110;
20'b01001001000110101111: color_data = 12'b111011101110;
20'b01001001000110110000: color_data = 12'b111011101110;
20'b01001001000110111101: color_data = 12'b111011101110;
20'b01001001000110111110: color_data = 12'b111011101110;
20'b01001001000110111111: color_data = 12'b111011101110;
20'b01001001000111000000: color_data = 12'b111011101110;
20'b01001001000111000001: color_data = 12'b111011101110;
20'b01001001000111000010: color_data = 12'b111011101110;
20'b01001001000111000011: color_data = 12'b111011101110;
20'b01001001000111000100: color_data = 12'b111011101110;
20'b01001001000111000101: color_data = 12'b111011101110;
20'b01001001000111000110: color_data = 12'b111011101110;
20'b01001001000111001000: color_data = 12'b111011101110;
20'b01001001000111001001: color_data = 12'b111011101110;
20'b01001001000111001010: color_data = 12'b111011101110;
20'b01001001000111001011: color_data = 12'b111011101110;
20'b01001001000111001100: color_data = 12'b111011101110;
20'b01001001000111001101: color_data = 12'b111011101110;
20'b01001001000111001110: color_data = 12'b111011101110;
20'b01001001000111001111: color_data = 12'b111011101110;
20'b01001001000111010000: color_data = 12'b111011101110;
20'b01001001000111010001: color_data = 12'b111011101110;
20'b01001001000111010011: color_data = 12'b111011101110;
20'b01001001000111010100: color_data = 12'b111011101110;
20'b01001001000111010101: color_data = 12'b111011101110;
20'b01001001000111010110: color_data = 12'b111011101110;
20'b01001001000111010111: color_data = 12'b111011101110;
20'b01001001000111011000: color_data = 12'b111011101110;
20'b01001001000111011001: color_data = 12'b111011101110;
20'b01001001000111011010: color_data = 12'b111011101110;
20'b01001001000111011011: color_data = 12'b111011101110;
20'b01001001000111011100: color_data = 12'b111011101110;
20'b01001001010010010110: color_data = 12'b111011101110;
20'b01001001010010010111: color_data = 12'b111011101110;
20'b01001001010010011000: color_data = 12'b111011101110;
20'b01001001010010011001: color_data = 12'b111011101110;
20'b01001001010010011010: color_data = 12'b111011101110;
20'b01001001010010011011: color_data = 12'b111011101110;
20'b01001001010010011100: color_data = 12'b111011101110;
20'b01001001010010011101: color_data = 12'b111011101110;
20'b01001001010010011110: color_data = 12'b111011101110;
20'b01001001010010011111: color_data = 12'b111011101110;
20'b01001001010010100001: color_data = 12'b111011101110;
20'b01001001010010100010: color_data = 12'b111011101110;
20'b01001001010010100011: color_data = 12'b111011101110;
20'b01001001010010100100: color_data = 12'b111011101110;
20'b01001001010010100101: color_data = 12'b111011101110;
20'b01001001010010100110: color_data = 12'b111011101110;
20'b01001001010010100111: color_data = 12'b111011101110;
20'b01001001010010101000: color_data = 12'b111011101110;
20'b01001001010010101001: color_data = 12'b111011101110;
20'b01001001010010101010: color_data = 12'b111011101110;
20'b01001001010011001101: color_data = 12'b111011101110;
20'b01001001010011001110: color_data = 12'b111011101110;
20'b01001001010011001111: color_data = 12'b111011101110;
20'b01001001010011010000: color_data = 12'b111011101110;
20'b01001001010011010001: color_data = 12'b111011101110;
20'b01001001010011010010: color_data = 12'b111011101110;
20'b01001001010011010011: color_data = 12'b111011101110;
20'b01001001010011010100: color_data = 12'b111011101110;
20'b01001001010011010101: color_data = 12'b111011101110;
20'b01001001010011010110: color_data = 12'b111011101110;
20'b01001001010011011000: color_data = 12'b111011101110;
20'b01001001010011011001: color_data = 12'b111011101110;
20'b01001001010011011010: color_data = 12'b111011101110;
20'b01001001010011011011: color_data = 12'b111011101110;
20'b01001001010011011100: color_data = 12'b111011101110;
20'b01001001010011011101: color_data = 12'b111011101110;
20'b01001001010011011110: color_data = 12'b111011101110;
20'b01001001010011011111: color_data = 12'b111011101110;
20'b01001001010011100000: color_data = 12'b111011101110;
20'b01001001010011100001: color_data = 12'b111011101110;
20'b01001001010011101101: color_data = 12'b111011101110;
20'b01001001010011101110: color_data = 12'b111011101110;
20'b01001001010011101111: color_data = 12'b111011101110;
20'b01001001010011110000: color_data = 12'b111011101110;
20'b01001001010011110001: color_data = 12'b111011101110;
20'b01001001010011110010: color_data = 12'b111011101110;
20'b01001001010011110011: color_data = 12'b111011101110;
20'b01001001010011110100: color_data = 12'b111011101110;
20'b01001001010011110101: color_data = 12'b111011101110;
20'b01001001010011110110: color_data = 12'b111011101110;
20'b01001001010011111000: color_data = 12'b111011101110;
20'b01001001010011111001: color_data = 12'b111011101110;
20'b01001001010011111010: color_data = 12'b111011101110;
20'b01001001010011111011: color_data = 12'b111011101110;
20'b01001001010011111100: color_data = 12'b111011101110;
20'b01001001010011111101: color_data = 12'b111011101110;
20'b01001001010011111110: color_data = 12'b111011101110;
20'b01001001010011111111: color_data = 12'b111011101110;
20'b01001001010100000000: color_data = 12'b111011101110;
20'b01001001010100000001: color_data = 12'b111011101110;
20'b01001001010100100100: color_data = 12'b111011101110;
20'b01001001010100100101: color_data = 12'b111011101110;
20'b01001001010100100110: color_data = 12'b111011101110;
20'b01001001010100100111: color_data = 12'b111011101110;
20'b01001001010100101000: color_data = 12'b111011101110;
20'b01001001010100101001: color_data = 12'b111011101110;
20'b01001001010100101010: color_data = 12'b111011101110;
20'b01001001010100101011: color_data = 12'b111011101110;
20'b01001001010100101100: color_data = 12'b111011101110;
20'b01001001010100101101: color_data = 12'b111011101110;
20'b01001001010100101111: color_data = 12'b111011101110;
20'b01001001010100110000: color_data = 12'b111011101110;
20'b01001001010100110001: color_data = 12'b111011101110;
20'b01001001010100110010: color_data = 12'b111011101110;
20'b01001001010100110011: color_data = 12'b111011101110;
20'b01001001010100110100: color_data = 12'b111011101110;
20'b01001001010100110101: color_data = 12'b111011101110;
20'b01001001010100110110: color_data = 12'b111011101110;
20'b01001001010100110111: color_data = 12'b111011101110;
20'b01001001010100111000: color_data = 12'b111011101110;
20'b01001001010101000100: color_data = 12'b111011101110;
20'b01001001010101000101: color_data = 12'b111011101110;
20'b01001001010101000110: color_data = 12'b111011101110;
20'b01001001010101000111: color_data = 12'b111011101110;
20'b01001001010101001000: color_data = 12'b111011101110;
20'b01001001010101001001: color_data = 12'b111011101110;
20'b01001001010101001010: color_data = 12'b111011101110;
20'b01001001010101001011: color_data = 12'b111011101110;
20'b01001001010101001100: color_data = 12'b111011101110;
20'b01001001010101001101: color_data = 12'b111011101110;
20'b01001001010101001111: color_data = 12'b111011101110;
20'b01001001010101010000: color_data = 12'b111011101110;
20'b01001001010101010001: color_data = 12'b111011101110;
20'b01001001010101010010: color_data = 12'b111011101110;
20'b01001001010101010011: color_data = 12'b111011101110;
20'b01001001010101010100: color_data = 12'b111011101110;
20'b01001001010101010101: color_data = 12'b111011101110;
20'b01001001010101010110: color_data = 12'b111011101110;
20'b01001001010101010111: color_data = 12'b111011101110;
20'b01001001010101011000: color_data = 12'b111011101110;
20'b01001001010101011010: color_data = 12'b111011101110;
20'b01001001010101011011: color_data = 12'b111011101110;
20'b01001001010101011100: color_data = 12'b111011101110;
20'b01001001010101011101: color_data = 12'b111011101110;
20'b01001001010101011110: color_data = 12'b111011101110;
20'b01001001010101011111: color_data = 12'b111011101110;
20'b01001001010101100000: color_data = 12'b111011101110;
20'b01001001010101100001: color_data = 12'b111011101110;
20'b01001001010101100010: color_data = 12'b111011101110;
20'b01001001010101100011: color_data = 12'b111011101110;
20'b01001001010101100101: color_data = 12'b111011101110;
20'b01001001010101100110: color_data = 12'b111011101110;
20'b01001001010101100111: color_data = 12'b111011101110;
20'b01001001010101101000: color_data = 12'b111011101110;
20'b01001001010101101001: color_data = 12'b111011101110;
20'b01001001010101101010: color_data = 12'b111011101110;
20'b01001001010101101011: color_data = 12'b111011101110;
20'b01001001010101101100: color_data = 12'b111011101110;
20'b01001001010101101101: color_data = 12'b111011101110;
20'b01001001010101101110: color_data = 12'b111011101110;
20'b01001001010101110000: color_data = 12'b111011101110;
20'b01001001010101110001: color_data = 12'b111011101110;
20'b01001001010101110010: color_data = 12'b111011101110;
20'b01001001010101110011: color_data = 12'b111011101110;
20'b01001001010101110100: color_data = 12'b111011101110;
20'b01001001010101110101: color_data = 12'b111011101110;
20'b01001001010101110110: color_data = 12'b111011101110;
20'b01001001010101110111: color_data = 12'b111011101110;
20'b01001001010101111000: color_data = 12'b111011101110;
20'b01001001010101111001: color_data = 12'b111011101110;
20'b01001001010110011100: color_data = 12'b111011101110;
20'b01001001010110011101: color_data = 12'b111011101110;
20'b01001001010110011110: color_data = 12'b111011101110;
20'b01001001010110011111: color_data = 12'b111011101110;
20'b01001001010110100000: color_data = 12'b111011101110;
20'b01001001010110100001: color_data = 12'b111011101110;
20'b01001001010110100010: color_data = 12'b111011101110;
20'b01001001010110100011: color_data = 12'b111011101110;
20'b01001001010110100100: color_data = 12'b111011101110;
20'b01001001010110100101: color_data = 12'b111011101110;
20'b01001001010110100111: color_data = 12'b111011101110;
20'b01001001010110101000: color_data = 12'b111011101110;
20'b01001001010110101001: color_data = 12'b111011101110;
20'b01001001010110101010: color_data = 12'b111011101110;
20'b01001001010110101011: color_data = 12'b111011101110;
20'b01001001010110101100: color_data = 12'b111011101110;
20'b01001001010110101101: color_data = 12'b111011101110;
20'b01001001010110101110: color_data = 12'b111011101110;
20'b01001001010110101111: color_data = 12'b111011101110;
20'b01001001010110110000: color_data = 12'b111011101110;
20'b01001001010110111101: color_data = 12'b111011101110;
20'b01001001010110111110: color_data = 12'b111011101110;
20'b01001001010110111111: color_data = 12'b111011101110;
20'b01001001010111000000: color_data = 12'b111011101110;
20'b01001001010111000001: color_data = 12'b111011101110;
20'b01001001010111000010: color_data = 12'b111011101110;
20'b01001001010111000011: color_data = 12'b111011101110;
20'b01001001010111000100: color_data = 12'b111011101110;
20'b01001001010111000101: color_data = 12'b111011101110;
20'b01001001010111000110: color_data = 12'b111011101110;
20'b01001001010111001000: color_data = 12'b111011101110;
20'b01001001010111001001: color_data = 12'b111011101110;
20'b01001001010111001010: color_data = 12'b111011101110;
20'b01001001010111001011: color_data = 12'b111011101110;
20'b01001001010111001100: color_data = 12'b111011101110;
20'b01001001010111001101: color_data = 12'b111011101110;
20'b01001001010111001110: color_data = 12'b111011101110;
20'b01001001010111001111: color_data = 12'b111011101110;
20'b01001001010111010000: color_data = 12'b111011101110;
20'b01001001010111010001: color_data = 12'b111011101110;
20'b01001001010111010011: color_data = 12'b111011101110;
20'b01001001010111010100: color_data = 12'b111011101110;
20'b01001001010111010101: color_data = 12'b111011101110;
20'b01001001010111010110: color_data = 12'b111011101110;
20'b01001001010111010111: color_data = 12'b111011101110;
20'b01001001010111011000: color_data = 12'b111011101110;
20'b01001001010111011001: color_data = 12'b111011101110;
20'b01001001010111011010: color_data = 12'b111011101110;
20'b01001001010111011011: color_data = 12'b111011101110;
20'b01001001010111011100: color_data = 12'b111011101110;
20'b01001001100010010110: color_data = 12'b111011101110;
20'b01001001100010010111: color_data = 12'b111011101110;
20'b01001001100010011000: color_data = 12'b111011101110;
20'b01001001100010011001: color_data = 12'b111011101110;
20'b01001001100010011010: color_data = 12'b111011101110;
20'b01001001100010011011: color_data = 12'b111011101110;
20'b01001001100010011100: color_data = 12'b111011101110;
20'b01001001100010011101: color_data = 12'b111011101110;
20'b01001001100010011110: color_data = 12'b111011101110;
20'b01001001100010011111: color_data = 12'b111011101110;
20'b01001001100010100001: color_data = 12'b111011101110;
20'b01001001100010100010: color_data = 12'b111011101110;
20'b01001001100010100011: color_data = 12'b111011101110;
20'b01001001100010100100: color_data = 12'b111011101110;
20'b01001001100010100101: color_data = 12'b111011101110;
20'b01001001100010100110: color_data = 12'b111011101110;
20'b01001001100010100111: color_data = 12'b111011101110;
20'b01001001100010101000: color_data = 12'b111011101110;
20'b01001001100010101001: color_data = 12'b111011101110;
20'b01001001100010101010: color_data = 12'b111011101110;
20'b01001001100011001101: color_data = 12'b111011101110;
20'b01001001100011001110: color_data = 12'b111011101110;
20'b01001001100011001111: color_data = 12'b111011101110;
20'b01001001100011010000: color_data = 12'b111011101110;
20'b01001001100011010001: color_data = 12'b111011101110;
20'b01001001100011010010: color_data = 12'b111011101110;
20'b01001001100011010011: color_data = 12'b111011101110;
20'b01001001100011010100: color_data = 12'b111011101110;
20'b01001001100011010101: color_data = 12'b111011101110;
20'b01001001100011010110: color_data = 12'b111011101110;
20'b01001001100011011000: color_data = 12'b111011101110;
20'b01001001100011011001: color_data = 12'b111011101110;
20'b01001001100011011010: color_data = 12'b111011101110;
20'b01001001100011011011: color_data = 12'b111011101110;
20'b01001001100011011100: color_data = 12'b111011101110;
20'b01001001100011011101: color_data = 12'b111011101110;
20'b01001001100011011110: color_data = 12'b111011101110;
20'b01001001100011011111: color_data = 12'b111011101110;
20'b01001001100011100000: color_data = 12'b111011101110;
20'b01001001100011100001: color_data = 12'b111011101110;
20'b01001001100011101101: color_data = 12'b111011101110;
20'b01001001100011101110: color_data = 12'b111011101110;
20'b01001001100011101111: color_data = 12'b111011101110;
20'b01001001100011110000: color_data = 12'b111011101110;
20'b01001001100011110001: color_data = 12'b111011101110;
20'b01001001100011110010: color_data = 12'b111011101110;
20'b01001001100011110011: color_data = 12'b111011101110;
20'b01001001100011110100: color_data = 12'b111011101110;
20'b01001001100011110101: color_data = 12'b111011101110;
20'b01001001100011110110: color_data = 12'b111011101110;
20'b01001001100011111000: color_data = 12'b111011101110;
20'b01001001100011111001: color_data = 12'b111011101110;
20'b01001001100011111010: color_data = 12'b111011101110;
20'b01001001100011111011: color_data = 12'b111011101110;
20'b01001001100011111100: color_data = 12'b111011101110;
20'b01001001100011111101: color_data = 12'b111011101110;
20'b01001001100011111110: color_data = 12'b111011101110;
20'b01001001100011111111: color_data = 12'b111011101110;
20'b01001001100100000000: color_data = 12'b111011101110;
20'b01001001100100000001: color_data = 12'b111011101110;
20'b01001001100100100100: color_data = 12'b111011101110;
20'b01001001100100100101: color_data = 12'b111011101110;
20'b01001001100100100110: color_data = 12'b111011101110;
20'b01001001100100100111: color_data = 12'b111011101110;
20'b01001001100100101000: color_data = 12'b111011101110;
20'b01001001100100101001: color_data = 12'b111011101110;
20'b01001001100100101010: color_data = 12'b111011101110;
20'b01001001100100101011: color_data = 12'b111011101110;
20'b01001001100100101100: color_data = 12'b111011101110;
20'b01001001100100101101: color_data = 12'b111011101110;
20'b01001001100100101111: color_data = 12'b111011101110;
20'b01001001100100110000: color_data = 12'b111011101110;
20'b01001001100100110001: color_data = 12'b111011101110;
20'b01001001100100110010: color_data = 12'b111011101110;
20'b01001001100100110011: color_data = 12'b111011101110;
20'b01001001100100110100: color_data = 12'b111011101110;
20'b01001001100100110101: color_data = 12'b111011101110;
20'b01001001100100110110: color_data = 12'b111011101110;
20'b01001001100100110111: color_data = 12'b111011101110;
20'b01001001100100111000: color_data = 12'b111011101110;
20'b01001001100101000100: color_data = 12'b111011101110;
20'b01001001100101000101: color_data = 12'b111011101110;
20'b01001001100101000110: color_data = 12'b111011101110;
20'b01001001100101000111: color_data = 12'b111011101110;
20'b01001001100101001000: color_data = 12'b111011101110;
20'b01001001100101001001: color_data = 12'b111011101110;
20'b01001001100101001010: color_data = 12'b111011101110;
20'b01001001100101001011: color_data = 12'b111011101110;
20'b01001001100101001100: color_data = 12'b111011101110;
20'b01001001100101001101: color_data = 12'b111011101110;
20'b01001001100101001111: color_data = 12'b111011101110;
20'b01001001100101010000: color_data = 12'b111011101110;
20'b01001001100101010001: color_data = 12'b111011101110;
20'b01001001100101010010: color_data = 12'b111011101110;
20'b01001001100101010011: color_data = 12'b111011101110;
20'b01001001100101010100: color_data = 12'b111011101110;
20'b01001001100101010101: color_data = 12'b111011101110;
20'b01001001100101010110: color_data = 12'b111011101110;
20'b01001001100101010111: color_data = 12'b111011101110;
20'b01001001100101011000: color_data = 12'b111011101110;
20'b01001001100101011010: color_data = 12'b111011101110;
20'b01001001100101011011: color_data = 12'b111011101110;
20'b01001001100101011100: color_data = 12'b111011101110;
20'b01001001100101011101: color_data = 12'b111011101110;
20'b01001001100101011110: color_data = 12'b111011101110;
20'b01001001100101011111: color_data = 12'b111011101110;
20'b01001001100101100000: color_data = 12'b111011101110;
20'b01001001100101100001: color_data = 12'b111011101110;
20'b01001001100101100010: color_data = 12'b111011101110;
20'b01001001100101100011: color_data = 12'b111011101110;
20'b01001001100101100101: color_data = 12'b111011101110;
20'b01001001100101100110: color_data = 12'b111011101110;
20'b01001001100101100111: color_data = 12'b111011101110;
20'b01001001100101101000: color_data = 12'b111011101110;
20'b01001001100101101001: color_data = 12'b111011101110;
20'b01001001100101101010: color_data = 12'b111011101110;
20'b01001001100101101011: color_data = 12'b111011101110;
20'b01001001100101101100: color_data = 12'b111011101110;
20'b01001001100101101101: color_data = 12'b111011101110;
20'b01001001100101101110: color_data = 12'b111011101110;
20'b01001001100101110000: color_data = 12'b111011101110;
20'b01001001100101110001: color_data = 12'b111011101110;
20'b01001001100101110010: color_data = 12'b111011101110;
20'b01001001100101110011: color_data = 12'b111011101110;
20'b01001001100101110100: color_data = 12'b111011101110;
20'b01001001100101110101: color_data = 12'b111011101110;
20'b01001001100101110110: color_data = 12'b111011101110;
20'b01001001100101110111: color_data = 12'b111011101110;
20'b01001001100101111000: color_data = 12'b111011101110;
20'b01001001100101111001: color_data = 12'b111011101110;
20'b01001001100110011100: color_data = 12'b111011101110;
20'b01001001100110011101: color_data = 12'b111011101110;
20'b01001001100110011110: color_data = 12'b111011101110;
20'b01001001100110011111: color_data = 12'b111011101110;
20'b01001001100110100000: color_data = 12'b111011101110;
20'b01001001100110100001: color_data = 12'b111011101110;
20'b01001001100110100010: color_data = 12'b111011101110;
20'b01001001100110100011: color_data = 12'b111011101110;
20'b01001001100110100100: color_data = 12'b111011101110;
20'b01001001100110100101: color_data = 12'b111011101110;
20'b01001001100110100111: color_data = 12'b111011101110;
20'b01001001100110101000: color_data = 12'b111011101110;
20'b01001001100110101001: color_data = 12'b111011101110;
20'b01001001100110101010: color_data = 12'b111011101110;
20'b01001001100110101011: color_data = 12'b111011101110;
20'b01001001100110101100: color_data = 12'b111011101110;
20'b01001001100110101101: color_data = 12'b111011101110;
20'b01001001100110101110: color_data = 12'b111011101110;
20'b01001001100110101111: color_data = 12'b111011101110;
20'b01001001100110110000: color_data = 12'b111011101110;
20'b01001001100110111101: color_data = 12'b111011101110;
20'b01001001100110111110: color_data = 12'b111011101110;
20'b01001001100110111111: color_data = 12'b111011101110;
20'b01001001100111000000: color_data = 12'b111011101110;
20'b01001001100111000001: color_data = 12'b111011101110;
20'b01001001100111000010: color_data = 12'b111011101110;
20'b01001001100111000011: color_data = 12'b111011101110;
20'b01001001100111000100: color_data = 12'b111011101110;
20'b01001001100111000101: color_data = 12'b111011101110;
20'b01001001100111000110: color_data = 12'b111011101110;
20'b01001001100111001000: color_data = 12'b111011101110;
20'b01001001100111001001: color_data = 12'b111011101110;
20'b01001001100111001010: color_data = 12'b111011101110;
20'b01001001100111001011: color_data = 12'b111011101110;
20'b01001001100111001100: color_data = 12'b111011101110;
20'b01001001100111001101: color_data = 12'b111011101110;
20'b01001001100111001110: color_data = 12'b111011101110;
20'b01001001100111001111: color_data = 12'b111011101110;
20'b01001001100111010000: color_data = 12'b111011101110;
20'b01001001100111010001: color_data = 12'b111011101110;
20'b01001001100111010011: color_data = 12'b111011101110;
20'b01001001100111010100: color_data = 12'b111011101110;
20'b01001001100111010101: color_data = 12'b111011101110;
20'b01001001100111010110: color_data = 12'b111011101110;
20'b01001001100111010111: color_data = 12'b111011101110;
20'b01001001100111011000: color_data = 12'b111011101110;
20'b01001001100111011001: color_data = 12'b111011101110;
20'b01001001100111011010: color_data = 12'b111011101110;
20'b01001001100111011011: color_data = 12'b111011101110;
20'b01001001100111011100: color_data = 12'b111011101110;
20'b01001001110010010110: color_data = 12'b111011101110;
20'b01001001110010010111: color_data = 12'b111011101110;
20'b01001001110010011000: color_data = 12'b111011101110;
20'b01001001110010011001: color_data = 12'b111011101110;
20'b01001001110010011010: color_data = 12'b111011101110;
20'b01001001110010011011: color_data = 12'b111011101110;
20'b01001001110010011100: color_data = 12'b111011101110;
20'b01001001110010011101: color_data = 12'b111011101110;
20'b01001001110010011110: color_data = 12'b111011101110;
20'b01001001110010011111: color_data = 12'b111011101110;
20'b01001001110010100001: color_data = 12'b111011101110;
20'b01001001110010100010: color_data = 12'b111011101110;
20'b01001001110010100011: color_data = 12'b111011101110;
20'b01001001110010100100: color_data = 12'b111011101110;
20'b01001001110010100101: color_data = 12'b111011101110;
20'b01001001110010100110: color_data = 12'b111011101110;
20'b01001001110010100111: color_data = 12'b111011101110;
20'b01001001110010101000: color_data = 12'b111011101110;
20'b01001001110010101001: color_data = 12'b111011101110;
20'b01001001110010101010: color_data = 12'b111011101110;
20'b01001001110011001101: color_data = 12'b111011101110;
20'b01001001110011001110: color_data = 12'b111011101110;
20'b01001001110011001111: color_data = 12'b111011101110;
20'b01001001110011010000: color_data = 12'b111011101110;
20'b01001001110011010001: color_data = 12'b111011101110;
20'b01001001110011010010: color_data = 12'b111011101110;
20'b01001001110011010011: color_data = 12'b111011101110;
20'b01001001110011010100: color_data = 12'b111011101110;
20'b01001001110011010101: color_data = 12'b111011101110;
20'b01001001110011010110: color_data = 12'b111011101110;
20'b01001001110011011000: color_data = 12'b111011101110;
20'b01001001110011011001: color_data = 12'b111011101110;
20'b01001001110011011010: color_data = 12'b111011101110;
20'b01001001110011011011: color_data = 12'b111011101110;
20'b01001001110011011100: color_data = 12'b111011101110;
20'b01001001110011011101: color_data = 12'b111011101110;
20'b01001001110011011110: color_data = 12'b111011101110;
20'b01001001110011011111: color_data = 12'b111011101110;
20'b01001001110011100000: color_data = 12'b111011101110;
20'b01001001110011100001: color_data = 12'b111011101110;
20'b01001001110011101101: color_data = 12'b111011101110;
20'b01001001110011101110: color_data = 12'b111011101110;
20'b01001001110011101111: color_data = 12'b111011101110;
20'b01001001110011110000: color_data = 12'b111011101110;
20'b01001001110011110001: color_data = 12'b111011101110;
20'b01001001110011110010: color_data = 12'b111011101110;
20'b01001001110011110011: color_data = 12'b111011101110;
20'b01001001110011110100: color_data = 12'b111011101110;
20'b01001001110011110101: color_data = 12'b111011101110;
20'b01001001110011110110: color_data = 12'b111011101110;
20'b01001001110011111000: color_data = 12'b111011101110;
20'b01001001110011111001: color_data = 12'b111011101110;
20'b01001001110011111010: color_data = 12'b111011101110;
20'b01001001110011111011: color_data = 12'b111011101110;
20'b01001001110011111100: color_data = 12'b111011101110;
20'b01001001110011111101: color_data = 12'b111011101110;
20'b01001001110011111110: color_data = 12'b111011101110;
20'b01001001110011111111: color_data = 12'b111011101110;
20'b01001001110100000000: color_data = 12'b111011101110;
20'b01001001110100000001: color_data = 12'b111011101110;
20'b01001001110100100100: color_data = 12'b111011101110;
20'b01001001110100100101: color_data = 12'b111011101110;
20'b01001001110100100110: color_data = 12'b111011101110;
20'b01001001110100100111: color_data = 12'b111011101110;
20'b01001001110100101000: color_data = 12'b111011101110;
20'b01001001110100101001: color_data = 12'b111011101110;
20'b01001001110100101010: color_data = 12'b111011101110;
20'b01001001110100101011: color_data = 12'b111011101110;
20'b01001001110100101100: color_data = 12'b111011101110;
20'b01001001110100101101: color_data = 12'b111011101110;
20'b01001001110100101111: color_data = 12'b111011101110;
20'b01001001110100110000: color_data = 12'b111011101110;
20'b01001001110100110001: color_data = 12'b111011101110;
20'b01001001110100110010: color_data = 12'b111011101110;
20'b01001001110100110011: color_data = 12'b111011101110;
20'b01001001110100110100: color_data = 12'b111011101110;
20'b01001001110100110101: color_data = 12'b111011101110;
20'b01001001110100110110: color_data = 12'b111011101110;
20'b01001001110100110111: color_data = 12'b111011101110;
20'b01001001110100111000: color_data = 12'b111011101110;
20'b01001001110101000100: color_data = 12'b111011101110;
20'b01001001110101000101: color_data = 12'b111011101110;
20'b01001001110101000110: color_data = 12'b111011101110;
20'b01001001110101000111: color_data = 12'b111011101110;
20'b01001001110101001000: color_data = 12'b111011101110;
20'b01001001110101001001: color_data = 12'b111011101110;
20'b01001001110101001010: color_data = 12'b111011101110;
20'b01001001110101001011: color_data = 12'b111011101110;
20'b01001001110101001100: color_data = 12'b111011101110;
20'b01001001110101001101: color_data = 12'b111011101110;
20'b01001001110101001111: color_data = 12'b111011101110;
20'b01001001110101010000: color_data = 12'b111011101110;
20'b01001001110101010001: color_data = 12'b111011101110;
20'b01001001110101010010: color_data = 12'b111011101110;
20'b01001001110101010011: color_data = 12'b111011101110;
20'b01001001110101010100: color_data = 12'b111011101110;
20'b01001001110101010101: color_data = 12'b111011101110;
20'b01001001110101010110: color_data = 12'b111011101110;
20'b01001001110101010111: color_data = 12'b111011101110;
20'b01001001110101011000: color_data = 12'b111011101110;
20'b01001001110101011010: color_data = 12'b111011101110;
20'b01001001110101011011: color_data = 12'b111011101110;
20'b01001001110101011100: color_data = 12'b111011101110;
20'b01001001110101011101: color_data = 12'b111011101110;
20'b01001001110101011110: color_data = 12'b111011101110;
20'b01001001110101011111: color_data = 12'b111011101110;
20'b01001001110101100000: color_data = 12'b111011101110;
20'b01001001110101100001: color_data = 12'b111011101110;
20'b01001001110101100010: color_data = 12'b111011101110;
20'b01001001110101100011: color_data = 12'b111011101110;
20'b01001001110101100101: color_data = 12'b111011101110;
20'b01001001110101100110: color_data = 12'b111011101110;
20'b01001001110101100111: color_data = 12'b111011101110;
20'b01001001110101101000: color_data = 12'b111011101110;
20'b01001001110101101001: color_data = 12'b111011101110;
20'b01001001110101101010: color_data = 12'b111011101110;
20'b01001001110101101011: color_data = 12'b111011101110;
20'b01001001110101101100: color_data = 12'b111011101110;
20'b01001001110101101101: color_data = 12'b111011101110;
20'b01001001110101101110: color_data = 12'b111011101110;
20'b01001001110101110000: color_data = 12'b111011101110;
20'b01001001110101110001: color_data = 12'b111011101110;
20'b01001001110101110010: color_data = 12'b111011101110;
20'b01001001110101110011: color_data = 12'b111011101110;
20'b01001001110101110100: color_data = 12'b111011101110;
20'b01001001110101110101: color_data = 12'b111011101110;
20'b01001001110101110110: color_data = 12'b111011101110;
20'b01001001110101110111: color_data = 12'b111011101110;
20'b01001001110101111000: color_data = 12'b111011101110;
20'b01001001110101111001: color_data = 12'b111011101110;
20'b01001001110110011100: color_data = 12'b111011101110;
20'b01001001110110011101: color_data = 12'b111011101110;
20'b01001001110110011110: color_data = 12'b111011101110;
20'b01001001110110011111: color_data = 12'b111011101110;
20'b01001001110110100000: color_data = 12'b111011101110;
20'b01001001110110100001: color_data = 12'b111011101110;
20'b01001001110110100010: color_data = 12'b111011101110;
20'b01001001110110100011: color_data = 12'b111011101110;
20'b01001001110110100100: color_data = 12'b111011101110;
20'b01001001110110100101: color_data = 12'b111011101110;
20'b01001001110110100111: color_data = 12'b111011101110;
20'b01001001110110101000: color_data = 12'b111011101110;
20'b01001001110110101001: color_data = 12'b111011101110;
20'b01001001110110101010: color_data = 12'b111011101110;
20'b01001001110110101011: color_data = 12'b111011101110;
20'b01001001110110101100: color_data = 12'b111011101110;
20'b01001001110110101101: color_data = 12'b111011101110;
20'b01001001110110101110: color_data = 12'b111011101110;
20'b01001001110110101111: color_data = 12'b111011101110;
20'b01001001110110110000: color_data = 12'b111011101110;
20'b01001001110110111101: color_data = 12'b111011101110;
20'b01001001110110111110: color_data = 12'b111011101110;
20'b01001001110110111111: color_data = 12'b111011101110;
20'b01001001110111000000: color_data = 12'b111011101110;
20'b01001001110111000001: color_data = 12'b111011101110;
20'b01001001110111000010: color_data = 12'b111011101110;
20'b01001001110111000011: color_data = 12'b111011101110;
20'b01001001110111000100: color_data = 12'b111011101110;
20'b01001001110111000101: color_data = 12'b111011101110;
20'b01001001110111000110: color_data = 12'b111011101110;
20'b01001001110111001000: color_data = 12'b111011101110;
20'b01001001110111001001: color_data = 12'b111011101110;
20'b01001001110111001010: color_data = 12'b111011101110;
20'b01001001110111001011: color_data = 12'b111011101110;
20'b01001001110111001100: color_data = 12'b111011101110;
20'b01001001110111001101: color_data = 12'b111011101110;
20'b01001001110111001110: color_data = 12'b111011101110;
20'b01001001110111001111: color_data = 12'b111011101110;
20'b01001001110111010000: color_data = 12'b111011101110;
20'b01001001110111010001: color_data = 12'b111011101110;
20'b01001001110111010011: color_data = 12'b111011101110;
20'b01001001110111010100: color_data = 12'b111011101110;
20'b01001001110111010101: color_data = 12'b111011101110;
20'b01001001110111010110: color_data = 12'b111011101110;
20'b01001001110111010111: color_data = 12'b111011101110;
20'b01001001110111011000: color_data = 12'b111011101110;
20'b01001001110111011001: color_data = 12'b111011101110;
20'b01001001110111011010: color_data = 12'b111011101110;
20'b01001001110111011011: color_data = 12'b111011101110;
20'b01001001110111011100: color_data = 12'b111011101110;
20'b01001010000010010110: color_data = 12'b111011101110;
20'b01001010000010010111: color_data = 12'b111011101110;
20'b01001010000010011000: color_data = 12'b111011101110;
20'b01001010000010011001: color_data = 12'b111011101110;
20'b01001010000010011010: color_data = 12'b111011101110;
20'b01001010000010011011: color_data = 12'b111011101110;
20'b01001010000010011100: color_data = 12'b111011101110;
20'b01001010000010011101: color_data = 12'b111011101110;
20'b01001010000010011110: color_data = 12'b111011101110;
20'b01001010000010011111: color_data = 12'b111011101110;
20'b01001010000010100001: color_data = 12'b111011101110;
20'b01001010000010100010: color_data = 12'b111011101110;
20'b01001010000010100011: color_data = 12'b111011101110;
20'b01001010000010100100: color_data = 12'b111011101110;
20'b01001010000010100101: color_data = 12'b111011101110;
20'b01001010000010100110: color_data = 12'b111011101110;
20'b01001010000010100111: color_data = 12'b111011101110;
20'b01001010000010101000: color_data = 12'b111011101110;
20'b01001010000010101001: color_data = 12'b111011101110;
20'b01001010000010101010: color_data = 12'b111011101110;
20'b01001010000011001101: color_data = 12'b111011101110;
20'b01001010000011001110: color_data = 12'b111011101110;
20'b01001010000011001111: color_data = 12'b111011101110;
20'b01001010000011010000: color_data = 12'b111011101110;
20'b01001010000011010001: color_data = 12'b111011101110;
20'b01001010000011010010: color_data = 12'b111011101110;
20'b01001010000011010011: color_data = 12'b111011101110;
20'b01001010000011010100: color_data = 12'b111011101110;
20'b01001010000011010101: color_data = 12'b111011101110;
20'b01001010000011010110: color_data = 12'b111011101110;
20'b01001010000011011000: color_data = 12'b111011101110;
20'b01001010000011011001: color_data = 12'b111011101110;
20'b01001010000011011010: color_data = 12'b111011101110;
20'b01001010000011011011: color_data = 12'b111011101110;
20'b01001010000011011100: color_data = 12'b111011101110;
20'b01001010000011011101: color_data = 12'b111011101110;
20'b01001010000011011110: color_data = 12'b111011101110;
20'b01001010000011011111: color_data = 12'b111011101110;
20'b01001010000011100000: color_data = 12'b111011101110;
20'b01001010000011100001: color_data = 12'b111011101110;
20'b01001010000011101101: color_data = 12'b111011101110;
20'b01001010000011101110: color_data = 12'b111011101110;
20'b01001010000011101111: color_data = 12'b111011101110;
20'b01001010000011110000: color_data = 12'b111011101110;
20'b01001010000011110001: color_data = 12'b111011101110;
20'b01001010000011110010: color_data = 12'b111011101110;
20'b01001010000011110011: color_data = 12'b111011101110;
20'b01001010000011110100: color_data = 12'b111011101110;
20'b01001010000011110101: color_data = 12'b111011101110;
20'b01001010000011110110: color_data = 12'b111011101110;
20'b01001010000011111000: color_data = 12'b111011101110;
20'b01001010000011111001: color_data = 12'b111011101110;
20'b01001010000011111010: color_data = 12'b111011101110;
20'b01001010000011111011: color_data = 12'b111011101110;
20'b01001010000011111100: color_data = 12'b111011101110;
20'b01001010000011111101: color_data = 12'b111011101110;
20'b01001010000011111110: color_data = 12'b111011101110;
20'b01001010000011111111: color_data = 12'b111011101110;
20'b01001010000100000000: color_data = 12'b111011101110;
20'b01001010000100000001: color_data = 12'b111011101110;
20'b01001010000100100100: color_data = 12'b111011101110;
20'b01001010000100100101: color_data = 12'b111011101110;
20'b01001010000100100110: color_data = 12'b111011101110;
20'b01001010000100100111: color_data = 12'b111011101110;
20'b01001010000100101000: color_data = 12'b111011101110;
20'b01001010000100101001: color_data = 12'b111011101110;
20'b01001010000100101010: color_data = 12'b111011101110;
20'b01001010000100101011: color_data = 12'b111011101110;
20'b01001010000100101100: color_data = 12'b111011101110;
20'b01001010000100101101: color_data = 12'b111011101110;
20'b01001010000100101111: color_data = 12'b111011101110;
20'b01001010000100110000: color_data = 12'b111011101110;
20'b01001010000100110001: color_data = 12'b111011101110;
20'b01001010000100110010: color_data = 12'b111011101110;
20'b01001010000100110011: color_data = 12'b111011101110;
20'b01001010000100110100: color_data = 12'b111011101110;
20'b01001010000100110101: color_data = 12'b111011101110;
20'b01001010000100110110: color_data = 12'b111011101110;
20'b01001010000100110111: color_data = 12'b111011101110;
20'b01001010000100111000: color_data = 12'b111011101110;
20'b01001010000101000100: color_data = 12'b111011101110;
20'b01001010000101000101: color_data = 12'b111011101110;
20'b01001010000101000110: color_data = 12'b111011101110;
20'b01001010000101000111: color_data = 12'b111011101110;
20'b01001010000101001000: color_data = 12'b111011101110;
20'b01001010000101001001: color_data = 12'b111011101110;
20'b01001010000101001010: color_data = 12'b111011101110;
20'b01001010000101001011: color_data = 12'b111011101110;
20'b01001010000101001100: color_data = 12'b111011101110;
20'b01001010000101001101: color_data = 12'b111011101110;
20'b01001010000101001111: color_data = 12'b111011101110;
20'b01001010000101010000: color_data = 12'b111011101110;
20'b01001010000101010001: color_data = 12'b111011101110;
20'b01001010000101010010: color_data = 12'b111011101110;
20'b01001010000101010011: color_data = 12'b111011101110;
20'b01001010000101010100: color_data = 12'b111011101110;
20'b01001010000101010101: color_data = 12'b111011101110;
20'b01001010000101010110: color_data = 12'b111011101110;
20'b01001010000101010111: color_data = 12'b111011101110;
20'b01001010000101011000: color_data = 12'b111011101110;
20'b01001010000101011010: color_data = 12'b111011101110;
20'b01001010000101011011: color_data = 12'b111011101110;
20'b01001010000101011100: color_data = 12'b111011101110;
20'b01001010000101011101: color_data = 12'b111011101110;
20'b01001010000101011110: color_data = 12'b111011101110;
20'b01001010000101011111: color_data = 12'b111011101110;
20'b01001010000101100000: color_data = 12'b111011101110;
20'b01001010000101100001: color_data = 12'b111011101110;
20'b01001010000101100010: color_data = 12'b111011101110;
20'b01001010000101100011: color_data = 12'b111011101110;
20'b01001010000101100101: color_data = 12'b111011101110;
20'b01001010000101100110: color_data = 12'b111011101110;
20'b01001010000101100111: color_data = 12'b111011101110;
20'b01001010000101101000: color_data = 12'b111011101110;
20'b01001010000101101001: color_data = 12'b111011101110;
20'b01001010000101101010: color_data = 12'b111011101110;
20'b01001010000101101011: color_data = 12'b111011101110;
20'b01001010000101101100: color_data = 12'b111011101110;
20'b01001010000101101101: color_data = 12'b111011101110;
20'b01001010000101101110: color_data = 12'b111011101110;
20'b01001010000101110000: color_data = 12'b111011101110;
20'b01001010000101110001: color_data = 12'b111011101110;
20'b01001010000101110010: color_data = 12'b111011101110;
20'b01001010000101110011: color_data = 12'b111011101110;
20'b01001010000101110100: color_data = 12'b111011101110;
20'b01001010000101110101: color_data = 12'b111011101110;
20'b01001010000101110110: color_data = 12'b111011101110;
20'b01001010000101110111: color_data = 12'b111011101110;
20'b01001010000101111000: color_data = 12'b111011101110;
20'b01001010000101111001: color_data = 12'b111011101110;
20'b01001010000110011100: color_data = 12'b111011101110;
20'b01001010000110011101: color_data = 12'b111011101110;
20'b01001010000110011110: color_data = 12'b111011101110;
20'b01001010000110011111: color_data = 12'b111011101110;
20'b01001010000110100000: color_data = 12'b111011101110;
20'b01001010000110100001: color_data = 12'b111011101110;
20'b01001010000110100010: color_data = 12'b111011101110;
20'b01001010000110100011: color_data = 12'b111011101110;
20'b01001010000110100100: color_data = 12'b111011101110;
20'b01001010000110100101: color_data = 12'b111011101110;
20'b01001010000110100111: color_data = 12'b111011101110;
20'b01001010000110101000: color_data = 12'b111011101110;
20'b01001010000110101001: color_data = 12'b111011101110;
20'b01001010000110101010: color_data = 12'b111011101110;
20'b01001010000110101011: color_data = 12'b111011101110;
20'b01001010000110101100: color_data = 12'b111011101110;
20'b01001010000110101101: color_data = 12'b111011101110;
20'b01001010000110101110: color_data = 12'b111011101110;
20'b01001010000110101111: color_data = 12'b111011101110;
20'b01001010000110110000: color_data = 12'b111011101110;
20'b01001010000110111101: color_data = 12'b111011101110;
20'b01001010000110111110: color_data = 12'b111011101110;
20'b01001010000110111111: color_data = 12'b111011101110;
20'b01001010000111000000: color_data = 12'b111011101110;
20'b01001010000111000001: color_data = 12'b111011101110;
20'b01001010000111000010: color_data = 12'b111011101110;
20'b01001010000111000011: color_data = 12'b111011101110;
20'b01001010000111000100: color_data = 12'b111011101110;
20'b01001010000111000101: color_data = 12'b111011101110;
20'b01001010000111000110: color_data = 12'b111011101110;
20'b01001010000111001000: color_data = 12'b111011101110;
20'b01001010000111001001: color_data = 12'b111011101110;
20'b01001010000111001010: color_data = 12'b111011101110;
20'b01001010000111001011: color_data = 12'b111011101110;
20'b01001010000111001100: color_data = 12'b111011101110;
20'b01001010000111001101: color_data = 12'b111011101110;
20'b01001010000111001110: color_data = 12'b111011101110;
20'b01001010000111001111: color_data = 12'b111011101110;
20'b01001010000111010000: color_data = 12'b111011101110;
20'b01001010000111010001: color_data = 12'b111011101110;
20'b01001010000111010011: color_data = 12'b111011101110;
20'b01001010000111010100: color_data = 12'b111011101110;
20'b01001010000111010101: color_data = 12'b111011101110;
20'b01001010000111010110: color_data = 12'b111011101110;
20'b01001010000111010111: color_data = 12'b111011101110;
20'b01001010000111011000: color_data = 12'b111011101110;
20'b01001010000111011001: color_data = 12'b111011101110;
20'b01001010000111011010: color_data = 12'b111011101110;
20'b01001010000111011011: color_data = 12'b111011101110;
20'b01001010000111011100: color_data = 12'b111011101110;
20'b01001010010010010110: color_data = 12'b111011101110;
20'b01001010010010010111: color_data = 12'b111011101110;
20'b01001010010010011000: color_data = 12'b111011101110;
20'b01001010010010011001: color_data = 12'b111011101110;
20'b01001010010010011010: color_data = 12'b111011101110;
20'b01001010010010011011: color_data = 12'b111011101110;
20'b01001010010010011100: color_data = 12'b111011101110;
20'b01001010010010011101: color_data = 12'b111011101110;
20'b01001010010010011110: color_data = 12'b111011101110;
20'b01001010010010011111: color_data = 12'b111011101110;
20'b01001010010010100001: color_data = 12'b111011101110;
20'b01001010010010100010: color_data = 12'b111011101110;
20'b01001010010010100011: color_data = 12'b111011101110;
20'b01001010010010100100: color_data = 12'b111011101110;
20'b01001010010010100101: color_data = 12'b111011101110;
20'b01001010010010100110: color_data = 12'b111011101110;
20'b01001010010010100111: color_data = 12'b111011101110;
20'b01001010010010101000: color_data = 12'b111011101110;
20'b01001010010010101001: color_data = 12'b111011101110;
20'b01001010010010101010: color_data = 12'b111011101110;
20'b01001010010011001101: color_data = 12'b111011101110;
20'b01001010010011001110: color_data = 12'b111011101110;
20'b01001010010011001111: color_data = 12'b111011101110;
20'b01001010010011010000: color_data = 12'b111011101110;
20'b01001010010011010001: color_data = 12'b111011101110;
20'b01001010010011010010: color_data = 12'b111011101110;
20'b01001010010011010011: color_data = 12'b111011101110;
20'b01001010010011010100: color_data = 12'b111011101110;
20'b01001010010011010101: color_data = 12'b111011101110;
20'b01001010010011010110: color_data = 12'b111011101110;
20'b01001010010011011000: color_data = 12'b111011101110;
20'b01001010010011011001: color_data = 12'b111011101110;
20'b01001010010011011010: color_data = 12'b111011101110;
20'b01001010010011011011: color_data = 12'b111011101110;
20'b01001010010011011100: color_data = 12'b111011101110;
20'b01001010010011011101: color_data = 12'b111011101110;
20'b01001010010011011110: color_data = 12'b111011101110;
20'b01001010010011011111: color_data = 12'b111011101110;
20'b01001010010011100000: color_data = 12'b111011101110;
20'b01001010010011100001: color_data = 12'b111011101110;
20'b01001010010011101101: color_data = 12'b111011101110;
20'b01001010010011101110: color_data = 12'b111011101110;
20'b01001010010011101111: color_data = 12'b111011101110;
20'b01001010010011110000: color_data = 12'b111011101110;
20'b01001010010011110001: color_data = 12'b111011101110;
20'b01001010010011110010: color_data = 12'b111011101110;
20'b01001010010011110011: color_data = 12'b111011101110;
20'b01001010010011110100: color_data = 12'b111011101110;
20'b01001010010011110101: color_data = 12'b111011101110;
20'b01001010010011110110: color_data = 12'b111011101110;
20'b01001010010011111000: color_data = 12'b111011101110;
20'b01001010010011111001: color_data = 12'b111011101110;
20'b01001010010011111010: color_data = 12'b111011101110;
20'b01001010010011111011: color_data = 12'b111011101110;
20'b01001010010011111100: color_data = 12'b111011101110;
20'b01001010010011111101: color_data = 12'b111011101110;
20'b01001010010011111110: color_data = 12'b111011101110;
20'b01001010010011111111: color_data = 12'b111011101110;
20'b01001010010100000000: color_data = 12'b111011101110;
20'b01001010010100000001: color_data = 12'b111011101110;
20'b01001010010100100100: color_data = 12'b111011101110;
20'b01001010010100100101: color_data = 12'b111011101110;
20'b01001010010100100110: color_data = 12'b111011101110;
20'b01001010010100100111: color_data = 12'b111011101110;
20'b01001010010100101000: color_data = 12'b111011101110;
20'b01001010010100101001: color_data = 12'b111011101110;
20'b01001010010100101010: color_data = 12'b111011101110;
20'b01001010010100101011: color_data = 12'b111011101110;
20'b01001010010100101100: color_data = 12'b111011101110;
20'b01001010010100101101: color_data = 12'b111011101110;
20'b01001010010100101111: color_data = 12'b111011101110;
20'b01001010010100110000: color_data = 12'b111011101110;
20'b01001010010100110001: color_data = 12'b111011101110;
20'b01001010010100110010: color_data = 12'b111011101110;
20'b01001010010100110011: color_data = 12'b111011101110;
20'b01001010010100110100: color_data = 12'b111011101110;
20'b01001010010100110101: color_data = 12'b111011101110;
20'b01001010010100110110: color_data = 12'b111011101110;
20'b01001010010100110111: color_data = 12'b111011101110;
20'b01001010010100111000: color_data = 12'b111011101110;
20'b01001010010101000100: color_data = 12'b111011101110;
20'b01001010010101000101: color_data = 12'b111011101110;
20'b01001010010101000110: color_data = 12'b111011101110;
20'b01001010010101000111: color_data = 12'b111011101110;
20'b01001010010101001000: color_data = 12'b111011101110;
20'b01001010010101001001: color_data = 12'b111011101110;
20'b01001010010101001010: color_data = 12'b111011101110;
20'b01001010010101001011: color_data = 12'b111011101110;
20'b01001010010101001100: color_data = 12'b111011101110;
20'b01001010010101001101: color_data = 12'b111011101110;
20'b01001010010101001111: color_data = 12'b111011101110;
20'b01001010010101010000: color_data = 12'b111011101110;
20'b01001010010101010001: color_data = 12'b111011101110;
20'b01001010010101010010: color_data = 12'b111011101110;
20'b01001010010101010011: color_data = 12'b111011101110;
20'b01001010010101010100: color_data = 12'b111011101110;
20'b01001010010101010101: color_data = 12'b111011101110;
20'b01001010010101010110: color_data = 12'b111011101110;
20'b01001010010101010111: color_data = 12'b111011101110;
20'b01001010010101011000: color_data = 12'b111011101110;
20'b01001010010101011010: color_data = 12'b111011101110;
20'b01001010010101011011: color_data = 12'b111011101110;
20'b01001010010101011100: color_data = 12'b111011101110;
20'b01001010010101011101: color_data = 12'b111011101110;
20'b01001010010101011110: color_data = 12'b111011101110;
20'b01001010010101011111: color_data = 12'b111011101110;
20'b01001010010101100000: color_data = 12'b111011101110;
20'b01001010010101100001: color_data = 12'b111011101110;
20'b01001010010101100010: color_data = 12'b111011101110;
20'b01001010010101100011: color_data = 12'b111011101110;
20'b01001010010101100101: color_data = 12'b111011101110;
20'b01001010010101100110: color_data = 12'b111011101110;
20'b01001010010101100111: color_data = 12'b111011101110;
20'b01001010010101101000: color_data = 12'b111011101110;
20'b01001010010101101001: color_data = 12'b111011101110;
20'b01001010010101101010: color_data = 12'b111011101110;
20'b01001010010101101011: color_data = 12'b111011101110;
20'b01001010010101101100: color_data = 12'b111011101110;
20'b01001010010101101101: color_data = 12'b111011101110;
20'b01001010010101101110: color_data = 12'b111011101110;
20'b01001010010101110000: color_data = 12'b111011101110;
20'b01001010010101110001: color_data = 12'b111011101110;
20'b01001010010101110010: color_data = 12'b111011101110;
20'b01001010010101110011: color_data = 12'b111011101110;
20'b01001010010101110100: color_data = 12'b111011101110;
20'b01001010010101110101: color_data = 12'b111011101110;
20'b01001010010101110110: color_data = 12'b111011101110;
20'b01001010010101110111: color_data = 12'b111011101110;
20'b01001010010101111000: color_data = 12'b111011101110;
20'b01001010010101111001: color_data = 12'b111011101110;
20'b01001010010110011100: color_data = 12'b111011101110;
20'b01001010010110011101: color_data = 12'b111011101110;
20'b01001010010110011110: color_data = 12'b111011101110;
20'b01001010010110011111: color_data = 12'b111011101110;
20'b01001010010110100000: color_data = 12'b111011101110;
20'b01001010010110100001: color_data = 12'b111011101110;
20'b01001010010110100010: color_data = 12'b111011101110;
20'b01001010010110100011: color_data = 12'b111011101110;
20'b01001010010110100100: color_data = 12'b111011101110;
20'b01001010010110100101: color_data = 12'b111011101110;
20'b01001010010110100111: color_data = 12'b111011101110;
20'b01001010010110101000: color_data = 12'b111011101110;
20'b01001010010110101001: color_data = 12'b111011101110;
20'b01001010010110101010: color_data = 12'b111011101110;
20'b01001010010110101011: color_data = 12'b111011101110;
20'b01001010010110101100: color_data = 12'b111011101110;
20'b01001010010110101101: color_data = 12'b111011101110;
20'b01001010010110101110: color_data = 12'b111011101110;
20'b01001010010110101111: color_data = 12'b111011101110;
20'b01001010010110110000: color_data = 12'b111011101110;
20'b01001010010110111101: color_data = 12'b111011101110;
20'b01001010010110111110: color_data = 12'b111011101110;
20'b01001010010110111111: color_data = 12'b111011101110;
20'b01001010010111000000: color_data = 12'b111011101110;
20'b01001010010111000001: color_data = 12'b111011101110;
20'b01001010010111000010: color_data = 12'b111011101110;
20'b01001010010111000011: color_data = 12'b111011101110;
20'b01001010010111000100: color_data = 12'b111011101110;
20'b01001010010111000101: color_data = 12'b111011101110;
20'b01001010010111000110: color_data = 12'b111011101110;
20'b01001010010111001000: color_data = 12'b111011101110;
20'b01001010010111001001: color_data = 12'b111011101110;
20'b01001010010111001010: color_data = 12'b111011101110;
20'b01001010010111001011: color_data = 12'b111011101110;
20'b01001010010111001100: color_data = 12'b111011101110;
20'b01001010010111001101: color_data = 12'b111011101110;
20'b01001010010111001110: color_data = 12'b111011101110;
20'b01001010010111001111: color_data = 12'b111011101110;
20'b01001010010111010000: color_data = 12'b111011101110;
20'b01001010010111010001: color_data = 12'b111011101110;
20'b01001010010111010011: color_data = 12'b111011101110;
20'b01001010010111010100: color_data = 12'b111011101110;
20'b01001010010111010101: color_data = 12'b111011101110;
20'b01001010010111010110: color_data = 12'b111011101110;
20'b01001010010111010111: color_data = 12'b111011101110;
20'b01001010010111011000: color_data = 12'b111011101110;
20'b01001010010111011001: color_data = 12'b111011101110;
20'b01001010010111011010: color_data = 12'b111011101110;
20'b01001010010111011011: color_data = 12'b111011101110;
20'b01001010010111011100: color_data = 12'b111011101110;
20'b01001010100010010110: color_data = 12'b111011101110;
20'b01001010100010010111: color_data = 12'b111011101110;
20'b01001010100010011000: color_data = 12'b111011101110;
20'b01001010100010011001: color_data = 12'b111011101110;
20'b01001010100010011010: color_data = 12'b111011101110;
20'b01001010100010011011: color_data = 12'b111011101110;
20'b01001010100010011100: color_data = 12'b111011101110;
20'b01001010100010011101: color_data = 12'b111011101110;
20'b01001010100010011110: color_data = 12'b111011101110;
20'b01001010100010011111: color_data = 12'b111011101110;
20'b01001010100010100001: color_data = 12'b111011101110;
20'b01001010100010100010: color_data = 12'b111011101110;
20'b01001010100010100011: color_data = 12'b111011101110;
20'b01001010100010100100: color_data = 12'b111011101110;
20'b01001010100010100101: color_data = 12'b111011101110;
20'b01001010100010100110: color_data = 12'b111011101110;
20'b01001010100010100111: color_data = 12'b111011101110;
20'b01001010100010101000: color_data = 12'b111011101110;
20'b01001010100010101001: color_data = 12'b111011101110;
20'b01001010100010101010: color_data = 12'b111011101110;
20'b01001010100011001101: color_data = 12'b111011101110;
20'b01001010100011001110: color_data = 12'b111011101110;
20'b01001010100011001111: color_data = 12'b111011101110;
20'b01001010100011010000: color_data = 12'b111011101110;
20'b01001010100011010001: color_data = 12'b111011101110;
20'b01001010100011010010: color_data = 12'b111011101110;
20'b01001010100011010011: color_data = 12'b111011101110;
20'b01001010100011010100: color_data = 12'b111011101110;
20'b01001010100011010101: color_data = 12'b111011101110;
20'b01001010100011010110: color_data = 12'b111011101110;
20'b01001010100011011000: color_data = 12'b111011101110;
20'b01001010100011011001: color_data = 12'b111011101110;
20'b01001010100011011010: color_data = 12'b111011101110;
20'b01001010100011011011: color_data = 12'b111011101110;
20'b01001010100011011100: color_data = 12'b111011101110;
20'b01001010100011011101: color_data = 12'b111011101110;
20'b01001010100011011110: color_data = 12'b111011101110;
20'b01001010100011011111: color_data = 12'b111011101110;
20'b01001010100011100000: color_data = 12'b111011101110;
20'b01001010100011100001: color_data = 12'b111011101110;
20'b01001010100011101101: color_data = 12'b111011101110;
20'b01001010100011101110: color_data = 12'b111011101110;
20'b01001010100011101111: color_data = 12'b111011101110;
20'b01001010100011110000: color_data = 12'b111011101110;
20'b01001010100011110001: color_data = 12'b111011101110;
20'b01001010100011110010: color_data = 12'b111011101110;
20'b01001010100011110011: color_data = 12'b111011101110;
20'b01001010100011110100: color_data = 12'b111011101110;
20'b01001010100011110101: color_data = 12'b111011101110;
20'b01001010100011110110: color_data = 12'b111011101110;
20'b01001010100011111000: color_data = 12'b111011101110;
20'b01001010100011111001: color_data = 12'b111011101110;
20'b01001010100011111010: color_data = 12'b111011101110;
20'b01001010100011111011: color_data = 12'b111011101110;
20'b01001010100011111100: color_data = 12'b111011101110;
20'b01001010100011111101: color_data = 12'b111011101110;
20'b01001010100011111110: color_data = 12'b111011101110;
20'b01001010100011111111: color_data = 12'b111011101110;
20'b01001010100100000000: color_data = 12'b111011101110;
20'b01001010100100000001: color_data = 12'b111011101110;
20'b01001010100100100100: color_data = 12'b111011101110;
20'b01001010100100100101: color_data = 12'b111011101110;
20'b01001010100100100110: color_data = 12'b111011101110;
20'b01001010100100100111: color_data = 12'b111011101110;
20'b01001010100100101000: color_data = 12'b111011101110;
20'b01001010100100101001: color_data = 12'b111011101110;
20'b01001010100100101010: color_data = 12'b111011101110;
20'b01001010100100101011: color_data = 12'b111011101110;
20'b01001010100100101100: color_data = 12'b111011101110;
20'b01001010100100101101: color_data = 12'b111011101110;
20'b01001010100100101111: color_data = 12'b111011101110;
20'b01001010100100110000: color_data = 12'b111011101110;
20'b01001010100100110001: color_data = 12'b111011101110;
20'b01001010100100110010: color_data = 12'b111011101110;
20'b01001010100100110011: color_data = 12'b111011101110;
20'b01001010100100110100: color_data = 12'b111011101110;
20'b01001010100100110101: color_data = 12'b111011101110;
20'b01001010100100110110: color_data = 12'b111011101110;
20'b01001010100100110111: color_data = 12'b111011101110;
20'b01001010100100111000: color_data = 12'b111011101110;
20'b01001010100101000100: color_data = 12'b111011101110;
20'b01001010100101000101: color_data = 12'b111011101110;
20'b01001010100101000110: color_data = 12'b111011101110;
20'b01001010100101000111: color_data = 12'b111011101110;
20'b01001010100101001000: color_data = 12'b111011101110;
20'b01001010100101001001: color_data = 12'b111011101110;
20'b01001010100101001010: color_data = 12'b111011101110;
20'b01001010100101001011: color_data = 12'b111011101110;
20'b01001010100101001100: color_data = 12'b111011101110;
20'b01001010100101001101: color_data = 12'b111011101110;
20'b01001010100101001111: color_data = 12'b111011101110;
20'b01001010100101010000: color_data = 12'b111011101110;
20'b01001010100101010001: color_data = 12'b111011101110;
20'b01001010100101010010: color_data = 12'b111011101110;
20'b01001010100101010011: color_data = 12'b111011101110;
20'b01001010100101010100: color_data = 12'b111011101110;
20'b01001010100101010101: color_data = 12'b111011101110;
20'b01001010100101010110: color_data = 12'b111011101110;
20'b01001010100101010111: color_data = 12'b111011101110;
20'b01001010100101011000: color_data = 12'b111011101110;
20'b01001010100101011010: color_data = 12'b111011101110;
20'b01001010100101011011: color_data = 12'b111011101110;
20'b01001010100101011100: color_data = 12'b111011101110;
20'b01001010100101011101: color_data = 12'b111011101110;
20'b01001010100101011110: color_data = 12'b111011101110;
20'b01001010100101011111: color_data = 12'b111011101110;
20'b01001010100101100000: color_data = 12'b111011101110;
20'b01001010100101100001: color_data = 12'b111011101110;
20'b01001010100101100010: color_data = 12'b111011101110;
20'b01001010100101100011: color_data = 12'b111011101110;
20'b01001010100101100101: color_data = 12'b111011101110;
20'b01001010100101100110: color_data = 12'b111011101110;
20'b01001010100101100111: color_data = 12'b111011101110;
20'b01001010100101101000: color_data = 12'b111011101110;
20'b01001010100101101001: color_data = 12'b111011101110;
20'b01001010100101101010: color_data = 12'b111011101110;
20'b01001010100101101011: color_data = 12'b111011101110;
20'b01001010100101101100: color_data = 12'b111011101110;
20'b01001010100101101101: color_data = 12'b111011101110;
20'b01001010100101101110: color_data = 12'b111011101110;
20'b01001010100101110000: color_data = 12'b111011101110;
20'b01001010100101110001: color_data = 12'b111011101110;
20'b01001010100101110010: color_data = 12'b111011101110;
20'b01001010100101110011: color_data = 12'b111011101110;
20'b01001010100101110100: color_data = 12'b111011101110;
20'b01001010100101110101: color_data = 12'b111011101110;
20'b01001010100101110110: color_data = 12'b111011101110;
20'b01001010100101110111: color_data = 12'b111011101110;
20'b01001010100101111000: color_data = 12'b111011101110;
20'b01001010100101111001: color_data = 12'b111011101110;
20'b01001010100110011100: color_data = 12'b111011101110;
20'b01001010100110011101: color_data = 12'b111011101110;
20'b01001010100110011110: color_data = 12'b111011101110;
20'b01001010100110011111: color_data = 12'b111011101110;
20'b01001010100110100000: color_data = 12'b111011101110;
20'b01001010100110100001: color_data = 12'b111011101110;
20'b01001010100110100010: color_data = 12'b111011101110;
20'b01001010100110100011: color_data = 12'b111011101110;
20'b01001010100110100100: color_data = 12'b111011101110;
20'b01001010100110100101: color_data = 12'b111011101110;
20'b01001010100110100111: color_data = 12'b111011101110;
20'b01001010100110101000: color_data = 12'b111011101110;
20'b01001010100110101001: color_data = 12'b111011101110;
20'b01001010100110101010: color_data = 12'b111011101110;
20'b01001010100110101011: color_data = 12'b111011101110;
20'b01001010100110101100: color_data = 12'b111011101110;
20'b01001010100110101101: color_data = 12'b111011101110;
20'b01001010100110101110: color_data = 12'b111011101110;
20'b01001010100110101111: color_data = 12'b111011101110;
20'b01001010100110110000: color_data = 12'b111011101110;
20'b01001010100110111101: color_data = 12'b111011101110;
20'b01001010100110111110: color_data = 12'b111011101110;
20'b01001010100110111111: color_data = 12'b111011101110;
20'b01001010100111000000: color_data = 12'b111011101110;
20'b01001010100111000001: color_data = 12'b111011101110;
20'b01001010100111000010: color_data = 12'b111011101110;
20'b01001010100111000011: color_data = 12'b111011101110;
20'b01001010100111000100: color_data = 12'b111011101110;
20'b01001010100111000101: color_data = 12'b111011101110;
20'b01001010100111000110: color_data = 12'b111011101110;
20'b01001010100111001000: color_data = 12'b111011101110;
20'b01001010100111001001: color_data = 12'b111011101110;
20'b01001010100111001010: color_data = 12'b111011101110;
20'b01001010100111001011: color_data = 12'b111011101110;
20'b01001010100111001100: color_data = 12'b111011101110;
20'b01001010100111001101: color_data = 12'b111011101110;
20'b01001010100111001110: color_data = 12'b111011101110;
20'b01001010100111001111: color_data = 12'b111011101110;
20'b01001010100111010000: color_data = 12'b111011101110;
20'b01001010100111010001: color_data = 12'b111011101110;
20'b01001010100111010011: color_data = 12'b111011101110;
20'b01001010100111010100: color_data = 12'b111011101110;
20'b01001010100111010101: color_data = 12'b111011101110;
20'b01001010100111010110: color_data = 12'b111011101110;
20'b01001010100111010111: color_data = 12'b111011101110;
20'b01001010100111011000: color_data = 12'b111011101110;
20'b01001010100111011001: color_data = 12'b111011101110;
20'b01001010100111011010: color_data = 12'b111011101110;
20'b01001010100111011011: color_data = 12'b111011101110;
20'b01001010100111011100: color_data = 12'b111011101110;
20'b01001011000010010110: color_data = 12'b111011101110;
20'b01001011000010010111: color_data = 12'b111011101110;
20'b01001011000010011000: color_data = 12'b111011101110;
20'b01001011000010011001: color_data = 12'b111011101110;
20'b01001011000010011010: color_data = 12'b111011101110;
20'b01001011000010011011: color_data = 12'b111011101110;
20'b01001011000010011100: color_data = 12'b111011101110;
20'b01001011000010011101: color_data = 12'b111011101110;
20'b01001011000010011110: color_data = 12'b111011101110;
20'b01001011000010011111: color_data = 12'b111011101110;
20'b01001011000010100001: color_data = 12'b111011101110;
20'b01001011000010100010: color_data = 12'b111011101110;
20'b01001011000010100011: color_data = 12'b111011101110;
20'b01001011000010100100: color_data = 12'b111011101110;
20'b01001011000010100101: color_data = 12'b111011101110;
20'b01001011000010100110: color_data = 12'b111011101110;
20'b01001011000010100111: color_data = 12'b111011101110;
20'b01001011000010101000: color_data = 12'b111011101110;
20'b01001011000010101001: color_data = 12'b111011101110;
20'b01001011000010101010: color_data = 12'b111011101110;
20'b01001011000011001101: color_data = 12'b111011101110;
20'b01001011000011001110: color_data = 12'b111011101110;
20'b01001011000011001111: color_data = 12'b111011101110;
20'b01001011000011010000: color_data = 12'b111011101110;
20'b01001011000011010001: color_data = 12'b111011101110;
20'b01001011000011010010: color_data = 12'b111011101110;
20'b01001011000011010011: color_data = 12'b111011101110;
20'b01001011000011010100: color_data = 12'b111011101110;
20'b01001011000011010101: color_data = 12'b111011101110;
20'b01001011000011010110: color_data = 12'b111011101110;
20'b01001011000011011000: color_data = 12'b111011101110;
20'b01001011000011011001: color_data = 12'b111011101110;
20'b01001011000011011010: color_data = 12'b111011101110;
20'b01001011000011011011: color_data = 12'b111011101110;
20'b01001011000011011100: color_data = 12'b111011101110;
20'b01001011000011011101: color_data = 12'b111011101110;
20'b01001011000011011110: color_data = 12'b111011101110;
20'b01001011000011011111: color_data = 12'b111011101110;
20'b01001011000011100000: color_data = 12'b111011101110;
20'b01001011000011100001: color_data = 12'b111011101110;
20'b01001011000011101101: color_data = 12'b111011101110;
20'b01001011000011101110: color_data = 12'b111011101110;
20'b01001011000011101111: color_data = 12'b111011101110;
20'b01001011000011110000: color_data = 12'b111011101110;
20'b01001011000011110001: color_data = 12'b111011101110;
20'b01001011000011110010: color_data = 12'b111011101110;
20'b01001011000011110011: color_data = 12'b111011101110;
20'b01001011000011110100: color_data = 12'b111011101110;
20'b01001011000011110101: color_data = 12'b111011101110;
20'b01001011000011110110: color_data = 12'b111011101110;
20'b01001011000011111000: color_data = 12'b111011101110;
20'b01001011000011111001: color_data = 12'b111011101110;
20'b01001011000011111010: color_data = 12'b111011101110;
20'b01001011000011111011: color_data = 12'b111011101110;
20'b01001011000011111100: color_data = 12'b111011101110;
20'b01001011000011111101: color_data = 12'b111011101110;
20'b01001011000011111110: color_data = 12'b111011101110;
20'b01001011000011111111: color_data = 12'b111011101110;
20'b01001011000100000000: color_data = 12'b111011101110;
20'b01001011000100000001: color_data = 12'b111011101110;
20'b01001011000100100100: color_data = 12'b111011101110;
20'b01001011000100100101: color_data = 12'b111011101110;
20'b01001011000100100110: color_data = 12'b111011101110;
20'b01001011000100100111: color_data = 12'b111011101110;
20'b01001011000100101000: color_data = 12'b111011101110;
20'b01001011000100101001: color_data = 12'b111011101110;
20'b01001011000100101010: color_data = 12'b111011101110;
20'b01001011000100101011: color_data = 12'b111011101110;
20'b01001011000100101100: color_data = 12'b111011101110;
20'b01001011000100101101: color_data = 12'b111011101110;
20'b01001011000100101111: color_data = 12'b111011101110;
20'b01001011000100110000: color_data = 12'b111011101110;
20'b01001011000100110001: color_data = 12'b111011101110;
20'b01001011000100110010: color_data = 12'b111011101110;
20'b01001011000100110011: color_data = 12'b111011101110;
20'b01001011000100110100: color_data = 12'b111011101110;
20'b01001011000100110101: color_data = 12'b111011101110;
20'b01001011000100110110: color_data = 12'b111011101110;
20'b01001011000100110111: color_data = 12'b111011101110;
20'b01001011000100111000: color_data = 12'b111011101110;
20'b01001011000101000100: color_data = 12'b111011101110;
20'b01001011000101000101: color_data = 12'b111011101110;
20'b01001011000101000110: color_data = 12'b111011101110;
20'b01001011000101000111: color_data = 12'b111011101110;
20'b01001011000101001000: color_data = 12'b111011101110;
20'b01001011000101001001: color_data = 12'b111011101110;
20'b01001011000101001010: color_data = 12'b111011101110;
20'b01001011000101001011: color_data = 12'b111011101110;
20'b01001011000101001100: color_data = 12'b111011101110;
20'b01001011000101001101: color_data = 12'b111011101110;
20'b01001011000101001111: color_data = 12'b111011101110;
20'b01001011000101010000: color_data = 12'b111011101110;
20'b01001011000101010001: color_data = 12'b111011101110;
20'b01001011000101010010: color_data = 12'b111011101110;
20'b01001011000101010011: color_data = 12'b111011101110;
20'b01001011000101010100: color_data = 12'b111011101110;
20'b01001011000101010101: color_data = 12'b111011101110;
20'b01001011000101010110: color_data = 12'b111011101110;
20'b01001011000101010111: color_data = 12'b111011101110;
20'b01001011000101011000: color_data = 12'b111011101110;
20'b01001011000110011100: color_data = 12'b111011101110;
20'b01001011000110011101: color_data = 12'b111011101110;
20'b01001011000110011110: color_data = 12'b111011101110;
20'b01001011000110011111: color_data = 12'b111011101110;
20'b01001011000110100000: color_data = 12'b111011101110;
20'b01001011000110100001: color_data = 12'b111011101110;
20'b01001011000110100010: color_data = 12'b111011101110;
20'b01001011000110100011: color_data = 12'b111011101110;
20'b01001011000110100100: color_data = 12'b111011101110;
20'b01001011000110100101: color_data = 12'b111011101110;
20'b01001011000110100111: color_data = 12'b111011101110;
20'b01001011000110101000: color_data = 12'b111011101110;
20'b01001011000110101001: color_data = 12'b111011101110;
20'b01001011000110101010: color_data = 12'b111011101110;
20'b01001011000110101011: color_data = 12'b111011101110;
20'b01001011000110101100: color_data = 12'b111011101110;
20'b01001011000110101101: color_data = 12'b111011101110;
20'b01001011000110101110: color_data = 12'b111011101110;
20'b01001011000110101111: color_data = 12'b111011101110;
20'b01001011000110110000: color_data = 12'b111011101110;
20'b01001011000110110010: color_data = 12'b111011101110;
20'b01001011000110110011: color_data = 12'b111011101110;
20'b01001011000110110100: color_data = 12'b111011101110;
20'b01001011000110110101: color_data = 12'b111011101110;
20'b01001011000110110110: color_data = 12'b111011101110;
20'b01001011000110110111: color_data = 12'b111011101110;
20'b01001011000110111000: color_data = 12'b111011101110;
20'b01001011000110111001: color_data = 12'b111011101110;
20'b01001011000110111010: color_data = 12'b111011101110;
20'b01001011000110111011: color_data = 12'b111011101110;
20'b01001011000110111101: color_data = 12'b111011101110;
20'b01001011000110111110: color_data = 12'b111011101110;
20'b01001011000110111111: color_data = 12'b111011101110;
20'b01001011000111000000: color_data = 12'b111011101110;
20'b01001011000111000001: color_data = 12'b111011101110;
20'b01001011000111000010: color_data = 12'b111011101110;
20'b01001011000111000011: color_data = 12'b111011101110;
20'b01001011000111000100: color_data = 12'b111011101110;
20'b01001011000111000101: color_data = 12'b111011101110;
20'b01001011000111000110: color_data = 12'b111011101110;
20'b01001011010010010110: color_data = 12'b111011101110;
20'b01001011010010010111: color_data = 12'b111011101110;
20'b01001011010010011000: color_data = 12'b111011101110;
20'b01001011010010011001: color_data = 12'b111011101110;
20'b01001011010010011010: color_data = 12'b111011101110;
20'b01001011010010011011: color_data = 12'b111011101110;
20'b01001011010010011100: color_data = 12'b111011101110;
20'b01001011010010011101: color_data = 12'b111011101110;
20'b01001011010010011110: color_data = 12'b111011101110;
20'b01001011010010011111: color_data = 12'b111011101110;
20'b01001011010010100001: color_data = 12'b111011101110;
20'b01001011010010100010: color_data = 12'b111011101110;
20'b01001011010010100011: color_data = 12'b111011101110;
20'b01001011010010100100: color_data = 12'b111011101110;
20'b01001011010010100101: color_data = 12'b111011101110;
20'b01001011010010100110: color_data = 12'b111011101110;
20'b01001011010010100111: color_data = 12'b111011101110;
20'b01001011010010101000: color_data = 12'b111011101110;
20'b01001011010010101001: color_data = 12'b111011101110;
20'b01001011010010101010: color_data = 12'b111011101110;
20'b01001011010011001101: color_data = 12'b111011101110;
20'b01001011010011001110: color_data = 12'b111011101110;
20'b01001011010011001111: color_data = 12'b111011101110;
20'b01001011010011010000: color_data = 12'b111011101110;
20'b01001011010011010001: color_data = 12'b111011101110;
20'b01001011010011010010: color_data = 12'b111011101110;
20'b01001011010011010011: color_data = 12'b111011101110;
20'b01001011010011010100: color_data = 12'b111011101110;
20'b01001011010011010101: color_data = 12'b111011101110;
20'b01001011010011010110: color_data = 12'b111011101110;
20'b01001011010011011000: color_data = 12'b111011101110;
20'b01001011010011011001: color_data = 12'b111011101110;
20'b01001011010011011010: color_data = 12'b111011101110;
20'b01001011010011011011: color_data = 12'b111011101110;
20'b01001011010011011100: color_data = 12'b111011101110;
20'b01001011010011011101: color_data = 12'b111011101110;
20'b01001011010011011110: color_data = 12'b111011101110;
20'b01001011010011011111: color_data = 12'b111011101110;
20'b01001011010011100000: color_data = 12'b111011101110;
20'b01001011010011100001: color_data = 12'b111011101110;
20'b01001011010011101101: color_data = 12'b111011101110;
20'b01001011010011101110: color_data = 12'b111011101110;
20'b01001011010011101111: color_data = 12'b111011101110;
20'b01001011010011110000: color_data = 12'b111011101110;
20'b01001011010011110001: color_data = 12'b111011101110;
20'b01001011010011110010: color_data = 12'b111011101110;
20'b01001011010011110011: color_data = 12'b111011101110;
20'b01001011010011110100: color_data = 12'b111011101110;
20'b01001011010011110101: color_data = 12'b111011101110;
20'b01001011010011110110: color_data = 12'b111011101110;
20'b01001011010011111000: color_data = 12'b111011101110;
20'b01001011010011111001: color_data = 12'b111011101110;
20'b01001011010011111010: color_data = 12'b111011101110;
20'b01001011010011111011: color_data = 12'b111011101110;
20'b01001011010011111100: color_data = 12'b111011101110;
20'b01001011010011111101: color_data = 12'b111011101110;
20'b01001011010011111110: color_data = 12'b111011101110;
20'b01001011010011111111: color_data = 12'b111011101110;
20'b01001011010100000000: color_data = 12'b111011101110;
20'b01001011010100000001: color_data = 12'b111011101110;
20'b01001011010100100100: color_data = 12'b111011101110;
20'b01001011010100100101: color_data = 12'b111011101110;
20'b01001011010100100110: color_data = 12'b111011101110;
20'b01001011010100100111: color_data = 12'b111011101110;
20'b01001011010100101000: color_data = 12'b111011101110;
20'b01001011010100101001: color_data = 12'b111011101110;
20'b01001011010100101010: color_data = 12'b111011101110;
20'b01001011010100101011: color_data = 12'b111011101110;
20'b01001011010100101100: color_data = 12'b111011101110;
20'b01001011010100101101: color_data = 12'b111011101110;
20'b01001011010100101111: color_data = 12'b111011101110;
20'b01001011010100110000: color_data = 12'b111011101110;
20'b01001011010100110001: color_data = 12'b111011101110;
20'b01001011010100110010: color_data = 12'b111011101110;
20'b01001011010100110011: color_data = 12'b111011101110;
20'b01001011010100110100: color_data = 12'b111011101110;
20'b01001011010100110101: color_data = 12'b111011101110;
20'b01001011010100110110: color_data = 12'b111011101110;
20'b01001011010100110111: color_data = 12'b111011101110;
20'b01001011010100111000: color_data = 12'b111011101110;
20'b01001011010101000100: color_data = 12'b111011101110;
20'b01001011010101000101: color_data = 12'b111011101110;
20'b01001011010101000110: color_data = 12'b111011101110;
20'b01001011010101000111: color_data = 12'b111011101110;
20'b01001011010101001000: color_data = 12'b111011101110;
20'b01001011010101001001: color_data = 12'b111011101110;
20'b01001011010101001010: color_data = 12'b111011101110;
20'b01001011010101001011: color_data = 12'b111011101110;
20'b01001011010101001100: color_data = 12'b111011101110;
20'b01001011010101001101: color_data = 12'b111011101110;
20'b01001011010101001111: color_data = 12'b111011101110;
20'b01001011010101010000: color_data = 12'b111011101110;
20'b01001011010101010001: color_data = 12'b111011101110;
20'b01001011010101010010: color_data = 12'b111011101110;
20'b01001011010101010011: color_data = 12'b111011101110;
20'b01001011010101010100: color_data = 12'b111011101110;
20'b01001011010101010101: color_data = 12'b111011101110;
20'b01001011010101010110: color_data = 12'b111011101110;
20'b01001011010101010111: color_data = 12'b111011101110;
20'b01001011010101011000: color_data = 12'b111011101110;
20'b01001011010110011100: color_data = 12'b111011101110;
20'b01001011010110011101: color_data = 12'b111011101110;
20'b01001011010110011110: color_data = 12'b111011101110;
20'b01001011010110011111: color_data = 12'b111011101110;
20'b01001011010110100000: color_data = 12'b111011101110;
20'b01001011010110100001: color_data = 12'b111011101110;
20'b01001011010110100010: color_data = 12'b111011101110;
20'b01001011010110100011: color_data = 12'b111011101110;
20'b01001011010110100100: color_data = 12'b111011101110;
20'b01001011010110100101: color_data = 12'b111011101110;
20'b01001011010110100111: color_data = 12'b111011101110;
20'b01001011010110101000: color_data = 12'b111011101110;
20'b01001011010110101001: color_data = 12'b111011101110;
20'b01001011010110101010: color_data = 12'b111011101110;
20'b01001011010110101011: color_data = 12'b111011101110;
20'b01001011010110101100: color_data = 12'b111011101110;
20'b01001011010110101101: color_data = 12'b111011101110;
20'b01001011010110101110: color_data = 12'b111011101110;
20'b01001011010110101111: color_data = 12'b111011101110;
20'b01001011010110110000: color_data = 12'b111011101110;
20'b01001011010110110010: color_data = 12'b111011101110;
20'b01001011010110110011: color_data = 12'b111011101110;
20'b01001011010110110100: color_data = 12'b111011101110;
20'b01001011010110110101: color_data = 12'b111011101110;
20'b01001011010110110110: color_data = 12'b111011101110;
20'b01001011010110110111: color_data = 12'b111011101110;
20'b01001011010110111000: color_data = 12'b111011101110;
20'b01001011010110111001: color_data = 12'b111011101110;
20'b01001011010110111010: color_data = 12'b111011101110;
20'b01001011010110111011: color_data = 12'b111011101110;
20'b01001011010110111101: color_data = 12'b111011101110;
20'b01001011010110111110: color_data = 12'b111011101110;
20'b01001011010110111111: color_data = 12'b111011101110;
20'b01001011010111000000: color_data = 12'b111011101110;
20'b01001011010111000001: color_data = 12'b111011101110;
20'b01001011010111000010: color_data = 12'b111011101110;
20'b01001011010111000011: color_data = 12'b111011101110;
20'b01001011010111000100: color_data = 12'b111011101110;
20'b01001011010111000101: color_data = 12'b111011101110;
20'b01001011010111000110: color_data = 12'b111011101110;
20'b01001011100010010110: color_data = 12'b111011101110;
20'b01001011100010010111: color_data = 12'b111011101110;
20'b01001011100010011000: color_data = 12'b111011101110;
20'b01001011100010011001: color_data = 12'b111011101110;
20'b01001011100010011010: color_data = 12'b111011101110;
20'b01001011100010011011: color_data = 12'b111011101110;
20'b01001011100010011100: color_data = 12'b111011101110;
20'b01001011100010011101: color_data = 12'b111011101110;
20'b01001011100010011110: color_data = 12'b111011101110;
20'b01001011100010011111: color_data = 12'b111011101110;
20'b01001011100010100001: color_data = 12'b111011101110;
20'b01001011100010100010: color_data = 12'b111011101110;
20'b01001011100010100011: color_data = 12'b111011101110;
20'b01001011100010100100: color_data = 12'b111011101110;
20'b01001011100010100101: color_data = 12'b111011101110;
20'b01001011100010100110: color_data = 12'b111011101110;
20'b01001011100010100111: color_data = 12'b111011101110;
20'b01001011100010101000: color_data = 12'b111011101110;
20'b01001011100010101001: color_data = 12'b111011101110;
20'b01001011100010101010: color_data = 12'b111011101110;
20'b01001011100011001101: color_data = 12'b111011101110;
20'b01001011100011001110: color_data = 12'b111011101110;
20'b01001011100011001111: color_data = 12'b111011101110;
20'b01001011100011010000: color_data = 12'b111011101110;
20'b01001011100011010001: color_data = 12'b111011101110;
20'b01001011100011010010: color_data = 12'b111011101110;
20'b01001011100011010011: color_data = 12'b111011101110;
20'b01001011100011010100: color_data = 12'b111011101110;
20'b01001011100011010101: color_data = 12'b111011101110;
20'b01001011100011010110: color_data = 12'b111011101110;
20'b01001011100011011000: color_data = 12'b111011101110;
20'b01001011100011011001: color_data = 12'b111011101110;
20'b01001011100011011010: color_data = 12'b111011101110;
20'b01001011100011011011: color_data = 12'b111011101110;
20'b01001011100011011100: color_data = 12'b111011101110;
20'b01001011100011011101: color_data = 12'b111011101110;
20'b01001011100011011110: color_data = 12'b111011101110;
20'b01001011100011011111: color_data = 12'b111011101110;
20'b01001011100011100000: color_data = 12'b111011101110;
20'b01001011100011100001: color_data = 12'b111011101110;
20'b01001011100011101101: color_data = 12'b111011101110;
20'b01001011100011101110: color_data = 12'b111011101110;
20'b01001011100011101111: color_data = 12'b111011101110;
20'b01001011100011110000: color_data = 12'b111011101110;
20'b01001011100011110001: color_data = 12'b111011101110;
20'b01001011100011110010: color_data = 12'b111011101110;
20'b01001011100011110011: color_data = 12'b111011101110;
20'b01001011100011110100: color_data = 12'b111011101110;
20'b01001011100011110101: color_data = 12'b111011101110;
20'b01001011100011110110: color_data = 12'b111011101110;
20'b01001011100011111000: color_data = 12'b111011101110;
20'b01001011100011111001: color_data = 12'b111011101110;
20'b01001011100011111010: color_data = 12'b111011101110;
20'b01001011100011111011: color_data = 12'b111011101110;
20'b01001011100011111100: color_data = 12'b111011101110;
20'b01001011100011111101: color_data = 12'b111011101110;
20'b01001011100011111110: color_data = 12'b111011101110;
20'b01001011100011111111: color_data = 12'b111011101110;
20'b01001011100100000000: color_data = 12'b111011101110;
20'b01001011100100000001: color_data = 12'b111011101110;
20'b01001011100100100100: color_data = 12'b111011101110;
20'b01001011100100100101: color_data = 12'b111011101110;
20'b01001011100100100110: color_data = 12'b111011101110;
20'b01001011100100100111: color_data = 12'b111011101110;
20'b01001011100100101000: color_data = 12'b111011101110;
20'b01001011100100101001: color_data = 12'b111011101110;
20'b01001011100100101010: color_data = 12'b111011101110;
20'b01001011100100101011: color_data = 12'b111011101110;
20'b01001011100100101100: color_data = 12'b111011101110;
20'b01001011100100101101: color_data = 12'b111011101110;
20'b01001011100100101111: color_data = 12'b111011101110;
20'b01001011100100110000: color_data = 12'b111011101110;
20'b01001011100100110001: color_data = 12'b111011101110;
20'b01001011100100110010: color_data = 12'b111011101110;
20'b01001011100100110011: color_data = 12'b111011101110;
20'b01001011100100110100: color_data = 12'b111011101110;
20'b01001011100100110101: color_data = 12'b111011101110;
20'b01001011100100110110: color_data = 12'b111011101110;
20'b01001011100100110111: color_data = 12'b111011101110;
20'b01001011100100111000: color_data = 12'b111011101110;
20'b01001011100101000100: color_data = 12'b111011101110;
20'b01001011100101000101: color_data = 12'b111011101110;
20'b01001011100101000110: color_data = 12'b111011101110;
20'b01001011100101000111: color_data = 12'b111011101110;
20'b01001011100101001000: color_data = 12'b111011101110;
20'b01001011100101001001: color_data = 12'b111011101110;
20'b01001011100101001010: color_data = 12'b111011101110;
20'b01001011100101001011: color_data = 12'b111011101110;
20'b01001011100101001100: color_data = 12'b111011101110;
20'b01001011100101001101: color_data = 12'b111011101110;
20'b01001011100101001111: color_data = 12'b111011101110;
20'b01001011100101010000: color_data = 12'b111011101110;
20'b01001011100101010001: color_data = 12'b111011101110;
20'b01001011100101010010: color_data = 12'b111011101110;
20'b01001011100101010011: color_data = 12'b111011101110;
20'b01001011100101010100: color_data = 12'b111011101110;
20'b01001011100101010101: color_data = 12'b111011101110;
20'b01001011100101010110: color_data = 12'b111011101110;
20'b01001011100101010111: color_data = 12'b111011101110;
20'b01001011100101011000: color_data = 12'b111011101110;
20'b01001011100110011100: color_data = 12'b111011101110;
20'b01001011100110011101: color_data = 12'b111011101110;
20'b01001011100110011110: color_data = 12'b111011101110;
20'b01001011100110011111: color_data = 12'b111011101110;
20'b01001011100110100000: color_data = 12'b111011101110;
20'b01001011100110100001: color_data = 12'b111011101110;
20'b01001011100110100010: color_data = 12'b111011101110;
20'b01001011100110100011: color_data = 12'b111011101110;
20'b01001011100110100100: color_data = 12'b111011101110;
20'b01001011100110100101: color_data = 12'b111011101110;
20'b01001011100110100111: color_data = 12'b111011101110;
20'b01001011100110101000: color_data = 12'b111011101110;
20'b01001011100110101001: color_data = 12'b111011101110;
20'b01001011100110101010: color_data = 12'b111011101110;
20'b01001011100110101011: color_data = 12'b111011101110;
20'b01001011100110101100: color_data = 12'b111011101110;
20'b01001011100110101101: color_data = 12'b111011101110;
20'b01001011100110101110: color_data = 12'b111011101110;
20'b01001011100110101111: color_data = 12'b111011101110;
20'b01001011100110110000: color_data = 12'b111011101110;
20'b01001011100110110010: color_data = 12'b111011101110;
20'b01001011100110110011: color_data = 12'b111011101110;
20'b01001011100110110100: color_data = 12'b111011101110;
20'b01001011100110110101: color_data = 12'b111011101110;
20'b01001011100110110110: color_data = 12'b111011101110;
20'b01001011100110110111: color_data = 12'b111011101110;
20'b01001011100110111000: color_data = 12'b111011101110;
20'b01001011100110111001: color_data = 12'b111011101110;
20'b01001011100110111010: color_data = 12'b111011101110;
20'b01001011100110111011: color_data = 12'b111011101110;
20'b01001011100110111101: color_data = 12'b111011101110;
20'b01001011100110111110: color_data = 12'b111011101110;
20'b01001011100110111111: color_data = 12'b111011101110;
20'b01001011100111000000: color_data = 12'b111011101110;
20'b01001011100111000001: color_data = 12'b111011101110;
20'b01001011100111000010: color_data = 12'b111011101110;
20'b01001011100111000011: color_data = 12'b111011101110;
20'b01001011100111000100: color_data = 12'b111011101110;
20'b01001011100111000101: color_data = 12'b111011101110;
20'b01001011100111000110: color_data = 12'b111011101110;
20'b01001011110010010110: color_data = 12'b111011101110;
20'b01001011110010010111: color_data = 12'b111011101110;
20'b01001011110010011000: color_data = 12'b111011101110;
20'b01001011110010011001: color_data = 12'b111011101110;
20'b01001011110010011010: color_data = 12'b111011101110;
20'b01001011110010011011: color_data = 12'b111011101110;
20'b01001011110010011100: color_data = 12'b111011101110;
20'b01001011110010011101: color_data = 12'b111011101110;
20'b01001011110010011110: color_data = 12'b111011101110;
20'b01001011110010011111: color_data = 12'b111011101110;
20'b01001011110010100001: color_data = 12'b111011101110;
20'b01001011110010100010: color_data = 12'b111011101110;
20'b01001011110010100011: color_data = 12'b111011101110;
20'b01001011110010100100: color_data = 12'b111011101110;
20'b01001011110010100101: color_data = 12'b111011101110;
20'b01001011110010100110: color_data = 12'b111011101110;
20'b01001011110010100111: color_data = 12'b111011101110;
20'b01001011110010101000: color_data = 12'b111011101110;
20'b01001011110010101001: color_data = 12'b111011101110;
20'b01001011110010101010: color_data = 12'b111011101110;
20'b01001011110011001101: color_data = 12'b111011101110;
20'b01001011110011001110: color_data = 12'b111011101110;
20'b01001011110011001111: color_data = 12'b111011101110;
20'b01001011110011010000: color_data = 12'b111011101110;
20'b01001011110011010001: color_data = 12'b111011101110;
20'b01001011110011010010: color_data = 12'b111011101110;
20'b01001011110011010011: color_data = 12'b111011101110;
20'b01001011110011010100: color_data = 12'b111011101110;
20'b01001011110011010101: color_data = 12'b111011101110;
20'b01001011110011010110: color_data = 12'b111011101110;
20'b01001011110011011000: color_data = 12'b111011101110;
20'b01001011110011011001: color_data = 12'b111011101110;
20'b01001011110011011010: color_data = 12'b111011101110;
20'b01001011110011011011: color_data = 12'b111011101110;
20'b01001011110011011100: color_data = 12'b111011101110;
20'b01001011110011011101: color_data = 12'b111011101110;
20'b01001011110011011110: color_data = 12'b111011101110;
20'b01001011110011011111: color_data = 12'b111011101110;
20'b01001011110011100000: color_data = 12'b111011101110;
20'b01001011110011100001: color_data = 12'b111011101110;
20'b01001011110011101101: color_data = 12'b111011101110;
20'b01001011110011101110: color_data = 12'b111011101110;
20'b01001011110011101111: color_data = 12'b111011101110;
20'b01001011110011110000: color_data = 12'b111011101110;
20'b01001011110011110001: color_data = 12'b111011101110;
20'b01001011110011110010: color_data = 12'b111011101110;
20'b01001011110011110011: color_data = 12'b111011101110;
20'b01001011110011110100: color_data = 12'b111011101110;
20'b01001011110011110101: color_data = 12'b111011101110;
20'b01001011110011110110: color_data = 12'b111011101110;
20'b01001011110011111000: color_data = 12'b111011101110;
20'b01001011110011111001: color_data = 12'b111011101110;
20'b01001011110011111010: color_data = 12'b111011101110;
20'b01001011110011111011: color_data = 12'b111011101110;
20'b01001011110011111100: color_data = 12'b111011101110;
20'b01001011110011111101: color_data = 12'b111011101110;
20'b01001011110011111110: color_data = 12'b111011101110;
20'b01001011110011111111: color_data = 12'b111011101110;
20'b01001011110100000000: color_data = 12'b111011101110;
20'b01001011110100000001: color_data = 12'b111011101110;
20'b01001011110100100100: color_data = 12'b111011101110;
20'b01001011110100100101: color_data = 12'b111011101110;
20'b01001011110100100110: color_data = 12'b111011101110;
20'b01001011110100100111: color_data = 12'b111011101110;
20'b01001011110100101000: color_data = 12'b111011101110;
20'b01001011110100101001: color_data = 12'b111011101110;
20'b01001011110100101010: color_data = 12'b111011101110;
20'b01001011110100101011: color_data = 12'b111011101110;
20'b01001011110100101100: color_data = 12'b111011101110;
20'b01001011110100101101: color_data = 12'b111011101110;
20'b01001011110100101111: color_data = 12'b111011101110;
20'b01001011110100110000: color_data = 12'b111011101110;
20'b01001011110100110001: color_data = 12'b111011101110;
20'b01001011110100110010: color_data = 12'b111011101110;
20'b01001011110100110011: color_data = 12'b111011101110;
20'b01001011110100110100: color_data = 12'b111011101110;
20'b01001011110100110101: color_data = 12'b111011101110;
20'b01001011110100110110: color_data = 12'b111011101110;
20'b01001011110100110111: color_data = 12'b111011101110;
20'b01001011110100111000: color_data = 12'b111011101110;
20'b01001011110101000100: color_data = 12'b111011101110;
20'b01001011110101000101: color_data = 12'b111011101110;
20'b01001011110101000110: color_data = 12'b111011101110;
20'b01001011110101000111: color_data = 12'b111011101110;
20'b01001011110101001000: color_data = 12'b111011101110;
20'b01001011110101001001: color_data = 12'b111011101110;
20'b01001011110101001010: color_data = 12'b111011101110;
20'b01001011110101001011: color_data = 12'b111011101110;
20'b01001011110101001100: color_data = 12'b111011101110;
20'b01001011110101001101: color_data = 12'b111011101110;
20'b01001011110101001111: color_data = 12'b111011101110;
20'b01001011110101010000: color_data = 12'b111011101110;
20'b01001011110101010001: color_data = 12'b111011101110;
20'b01001011110101010010: color_data = 12'b111011101110;
20'b01001011110101010011: color_data = 12'b111011101110;
20'b01001011110101010100: color_data = 12'b111011101110;
20'b01001011110101010101: color_data = 12'b111011101110;
20'b01001011110101010110: color_data = 12'b111011101110;
20'b01001011110101010111: color_data = 12'b111011101110;
20'b01001011110101011000: color_data = 12'b111011101110;
20'b01001011110110011100: color_data = 12'b111011101110;
20'b01001011110110011101: color_data = 12'b111011101110;
20'b01001011110110011110: color_data = 12'b111011101110;
20'b01001011110110011111: color_data = 12'b111011101110;
20'b01001011110110100000: color_data = 12'b111011101110;
20'b01001011110110100001: color_data = 12'b111011101110;
20'b01001011110110100010: color_data = 12'b111011101110;
20'b01001011110110100011: color_data = 12'b111011101110;
20'b01001011110110100100: color_data = 12'b111011101110;
20'b01001011110110100101: color_data = 12'b111011101110;
20'b01001011110110100111: color_data = 12'b111011101110;
20'b01001011110110101000: color_data = 12'b111011101110;
20'b01001011110110101001: color_data = 12'b111011101110;
20'b01001011110110101010: color_data = 12'b111011101110;
20'b01001011110110101011: color_data = 12'b111011101110;
20'b01001011110110101100: color_data = 12'b111011101110;
20'b01001011110110101101: color_data = 12'b111011101110;
20'b01001011110110101110: color_data = 12'b111011101110;
20'b01001011110110101111: color_data = 12'b111011101110;
20'b01001011110110110000: color_data = 12'b111011101110;
20'b01001011110110110010: color_data = 12'b111011101110;
20'b01001011110110110011: color_data = 12'b111011101110;
20'b01001011110110110100: color_data = 12'b111011101110;
20'b01001011110110110101: color_data = 12'b111011101110;
20'b01001011110110110110: color_data = 12'b111011101110;
20'b01001011110110110111: color_data = 12'b111011101110;
20'b01001011110110111000: color_data = 12'b111011101110;
20'b01001011110110111001: color_data = 12'b111011101110;
20'b01001011110110111010: color_data = 12'b111011101110;
20'b01001011110110111011: color_data = 12'b111011101110;
20'b01001011110110111101: color_data = 12'b111011101110;
20'b01001011110110111110: color_data = 12'b111011101110;
20'b01001011110110111111: color_data = 12'b111011101110;
20'b01001011110111000000: color_data = 12'b111011101110;
20'b01001011110111000001: color_data = 12'b111011101110;
20'b01001011110111000010: color_data = 12'b111011101110;
20'b01001011110111000011: color_data = 12'b111011101110;
20'b01001011110111000100: color_data = 12'b111011101110;
20'b01001011110111000101: color_data = 12'b111011101110;
20'b01001011110111000110: color_data = 12'b111011101110;
20'b01001100000010010110: color_data = 12'b111011101110;
20'b01001100000010010111: color_data = 12'b111011101110;
20'b01001100000010011000: color_data = 12'b111011101110;
20'b01001100000010011001: color_data = 12'b111011101110;
20'b01001100000010011010: color_data = 12'b111011101110;
20'b01001100000010011011: color_data = 12'b111011101110;
20'b01001100000010011100: color_data = 12'b111011101110;
20'b01001100000010011101: color_data = 12'b111011101110;
20'b01001100000010011110: color_data = 12'b111011101110;
20'b01001100000010011111: color_data = 12'b111011101110;
20'b01001100000010100001: color_data = 12'b111011101110;
20'b01001100000010100010: color_data = 12'b111011101110;
20'b01001100000010100011: color_data = 12'b111011101110;
20'b01001100000010100100: color_data = 12'b111011101110;
20'b01001100000010100101: color_data = 12'b111011101110;
20'b01001100000010100110: color_data = 12'b111011101110;
20'b01001100000010100111: color_data = 12'b111011101110;
20'b01001100000010101000: color_data = 12'b111011101110;
20'b01001100000010101001: color_data = 12'b111011101110;
20'b01001100000010101010: color_data = 12'b111011101110;
20'b01001100000011001101: color_data = 12'b111011101110;
20'b01001100000011001110: color_data = 12'b111011101110;
20'b01001100000011001111: color_data = 12'b111011101110;
20'b01001100000011010000: color_data = 12'b111011101110;
20'b01001100000011010001: color_data = 12'b111011101110;
20'b01001100000011010010: color_data = 12'b111011101110;
20'b01001100000011010011: color_data = 12'b111011101110;
20'b01001100000011010100: color_data = 12'b111011101110;
20'b01001100000011010101: color_data = 12'b111011101110;
20'b01001100000011010110: color_data = 12'b111011101110;
20'b01001100000011011000: color_data = 12'b111011101110;
20'b01001100000011011001: color_data = 12'b111011101110;
20'b01001100000011011010: color_data = 12'b111011101110;
20'b01001100000011011011: color_data = 12'b111011101110;
20'b01001100000011011100: color_data = 12'b111011101110;
20'b01001100000011011101: color_data = 12'b111011101110;
20'b01001100000011011110: color_data = 12'b111011101110;
20'b01001100000011011111: color_data = 12'b111011101110;
20'b01001100000011100000: color_data = 12'b111011101110;
20'b01001100000011100001: color_data = 12'b111011101110;
20'b01001100000011101101: color_data = 12'b111011101110;
20'b01001100000011101110: color_data = 12'b111011101110;
20'b01001100000011101111: color_data = 12'b111011101110;
20'b01001100000011110000: color_data = 12'b111011101110;
20'b01001100000011110001: color_data = 12'b111011101110;
20'b01001100000011110010: color_data = 12'b111011101110;
20'b01001100000011110011: color_data = 12'b111011101110;
20'b01001100000011110100: color_data = 12'b111011101110;
20'b01001100000011110101: color_data = 12'b111011101110;
20'b01001100000011110110: color_data = 12'b111011101110;
20'b01001100000011111000: color_data = 12'b111011101110;
20'b01001100000011111001: color_data = 12'b111011101110;
20'b01001100000011111010: color_data = 12'b111011101110;
20'b01001100000011111011: color_data = 12'b111011101110;
20'b01001100000011111100: color_data = 12'b111011101110;
20'b01001100000011111101: color_data = 12'b111011101110;
20'b01001100000011111110: color_data = 12'b111011101110;
20'b01001100000011111111: color_data = 12'b111011101110;
20'b01001100000100000000: color_data = 12'b111011101110;
20'b01001100000100000001: color_data = 12'b111011101110;
20'b01001100000100100100: color_data = 12'b111011101110;
20'b01001100000100100101: color_data = 12'b111011101110;
20'b01001100000100100110: color_data = 12'b111011101110;
20'b01001100000100100111: color_data = 12'b111011101110;
20'b01001100000100101000: color_data = 12'b111011101110;
20'b01001100000100101001: color_data = 12'b111011101110;
20'b01001100000100101010: color_data = 12'b111011101110;
20'b01001100000100101011: color_data = 12'b111011101110;
20'b01001100000100101100: color_data = 12'b111011101110;
20'b01001100000100101101: color_data = 12'b111011101110;
20'b01001100000100101111: color_data = 12'b111011101110;
20'b01001100000100110000: color_data = 12'b111011101110;
20'b01001100000100110001: color_data = 12'b111011101110;
20'b01001100000100110010: color_data = 12'b111011101110;
20'b01001100000100110011: color_data = 12'b111011101110;
20'b01001100000100110100: color_data = 12'b111011101110;
20'b01001100000100110101: color_data = 12'b111011101110;
20'b01001100000100110110: color_data = 12'b111011101110;
20'b01001100000100110111: color_data = 12'b111011101110;
20'b01001100000100111000: color_data = 12'b111011101110;
20'b01001100000101000100: color_data = 12'b111011101110;
20'b01001100000101000101: color_data = 12'b111011101110;
20'b01001100000101000110: color_data = 12'b111011101110;
20'b01001100000101000111: color_data = 12'b111011101110;
20'b01001100000101001000: color_data = 12'b111011101110;
20'b01001100000101001001: color_data = 12'b111011101110;
20'b01001100000101001010: color_data = 12'b111011101110;
20'b01001100000101001011: color_data = 12'b111011101110;
20'b01001100000101001100: color_data = 12'b111011101110;
20'b01001100000101001101: color_data = 12'b111011101110;
20'b01001100000101001111: color_data = 12'b111011101110;
20'b01001100000101010000: color_data = 12'b111011101110;
20'b01001100000101010001: color_data = 12'b111011101110;
20'b01001100000101010010: color_data = 12'b111011101110;
20'b01001100000101010011: color_data = 12'b111011101110;
20'b01001100000101010100: color_data = 12'b111011101110;
20'b01001100000101010101: color_data = 12'b111011101110;
20'b01001100000101010110: color_data = 12'b111011101110;
20'b01001100000101010111: color_data = 12'b111011101110;
20'b01001100000101011000: color_data = 12'b111011101110;
20'b01001100000110011100: color_data = 12'b111011101110;
20'b01001100000110011101: color_data = 12'b111011101110;
20'b01001100000110011110: color_data = 12'b111011101110;
20'b01001100000110011111: color_data = 12'b111011101110;
20'b01001100000110100000: color_data = 12'b111011101110;
20'b01001100000110100001: color_data = 12'b111011101110;
20'b01001100000110100010: color_data = 12'b111011101110;
20'b01001100000110100011: color_data = 12'b111011101110;
20'b01001100000110100100: color_data = 12'b111011101110;
20'b01001100000110100101: color_data = 12'b111011101110;
20'b01001100000110100111: color_data = 12'b111011101110;
20'b01001100000110101000: color_data = 12'b111011101110;
20'b01001100000110101001: color_data = 12'b111011101110;
20'b01001100000110101010: color_data = 12'b111011101110;
20'b01001100000110101011: color_data = 12'b111011101110;
20'b01001100000110101100: color_data = 12'b111011101110;
20'b01001100000110101101: color_data = 12'b111011101110;
20'b01001100000110101110: color_data = 12'b111011101110;
20'b01001100000110101111: color_data = 12'b111011101110;
20'b01001100000110110000: color_data = 12'b111011101110;
20'b01001100000110110010: color_data = 12'b111011101110;
20'b01001100000110110011: color_data = 12'b111011101110;
20'b01001100000110110100: color_data = 12'b111011101110;
20'b01001100000110110101: color_data = 12'b111011101110;
20'b01001100000110110110: color_data = 12'b111011101110;
20'b01001100000110110111: color_data = 12'b111011101110;
20'b01001100000110111000: color_data = 12'b111011101110;
20'b01001100000110111001: color_data = 12'b111011101110;
20'b01001100000110111010: color_data = 12'b111011101110;
20'b01001100000110111011: color_data = 12'b111011101110;
20'b01001100000110111101: color_data = 12'b111011101110;
20'b01001100000110111110: color_data = 12'b111011101110;
20'b01001100000110111111: color_data = 12'b111011101110;
20'b01001100000111000000: color_data = 12'b111011101110;
20'b01001100000111000001: color_data = 12'b111011101110;
20'b01001100000111000010: color_data = 12'b111011101110;
20'b01001100000111000011: color_data = 12'b111011101110;
20'b01001100000111000100: color_data = 12'b111011101110;
20'b01001100000111000101: color_data = 12'b111011101110;
20'b01001100000111000110: color_data = 12'b111011101110;
20'b01001100010010010110: color_data = 12'b111011101110;
20'b01001100010010010111: color_data = 12'b111011101110;
20'b01001100010010011000: color_data = 12'b111011101110;
20'b01001100010010011001: color_data = 12'b111011101110;
20'b01001100010010011010: color_data = 12'b111011101110;
20'b01001100010010011011: color_data = 12'b111011101110;
20'b01001100010010011100: color_data = 12'b111011101110;
20'b01001100010010011101: color_data = 12'b111011101110;
20'b01001100010010011110: color_data = 12'b111011101110;
20'b01001100010010011111: color_data = 12'b111011101110;
20'b01001100010010100001: color_data = 12'b111011101110;
20'b01001100010010100010: color_data = 12'b111011101110;
20'b01001100010010100011: color_data = 12'b111011101110;
20'b01001100010010100100: color_data = 12'b111011101110;
20'b01001100010010100101: color_data = 12'b111011101110;
20'b01001100010010100110: color_data = 12'b111011101110;
20'b01001100010010100111: color_data = 12'b111011101110;
20'b01001100010010101000: color_data = 12'b111011101110;
20'b01001100010010101001: color_data = 12'b111011101110;
20'b01001100010010101010: color_data = 12'b111011101110;
20'b01001100010011001101: color_data = 12'b111011101110;
20'b01001100010011001110: color_data = 12'b111011101110;
20'b01001100010011001111: color_data = 12'b111011101110;
20'b01001100010011010000: color_data = 12'b111011101110;
20'b01001100010011010001: color_data = 12'b111011101110;
20'b01001100010011010010: color_data = 12'b111011101110;
20'b01001100010011010011: color_data = 12'b111011101110;
20'b01001100010011010100: color_data = 12'b111011101110;
20'b01001100010011010101: color_data = 12'b111011101110;
20'b01001100010011010110: color_data = 12'b111011101110;
20'b01001100010011011000: color_data = 12'b111011101110;
20'b01001100010011011001: color_data = 12'b111011101110;
20'b01001100010011011010: color_data = 12'b111011101110;
20'b01001100010011011011: color_data = 12'b111011101110;
20'b01001100010011011100: color_data = 12'b111011101110;
20'b01001100010011011101: color_data = 12'b111011101110;
20'b01001100010011011110: color_data = 12'b111011101110;
20'b01001100010011011111: color_data = 12'b111011101110;
20'b01001100010011100000: color_data = 12'b111011101110;
20'b01001100010011100001: color_data = 12'b111011101110;
20'b01001100010011101101: color_data = 12'b111011101110;
20'b01001100010011101110: color_data = 12'b111011101110;
20'b01001100010011101111: color_data = 12'b111011101110;
20'b01001100010011110000: color_data = 12'b111011101110;
20'b01001100010011110001: color_data = 12'b111011101110;
20'b01001100010011110010: color_data = 12'b111011101110;
20'b01001100010011110011: color_data = 12'b111011101110;
20'b01001100010011110100: color_data = 12'b111011101110;
20'b01001100010011110101: color_data = 12'b111011101110;
20'b01001100010011110110: color_data = 12'b111011101110;
20'b01001100010011111000: color_data = 12'b111011101110;
20'b01001100010011111001: color_data = 12'b111011101110;
20'b01001100010011111010: color_data = 12'b111011101110;
20'b01001100010011111011: color_data = 12'b111011101110;
20'b01001100010011111100: color_data = 12'b111011101110;
20'b01001100010011111101: color_data = 12'b111011101110;
20'b01001100010011111110: color_data = 12'b111011101110;
20'b01001100010011111111: color_data = 12'b111011101110;
20'b01001100010100000000: color_data = 12'b111011101110;
20'b01001100010100000001: color_data = 12'b111011101110;
20'b01001100010100100100: color_data = 12'b111011101110;
20'b01001100010100100101: color_data = 12'b111011101110;
20'b01001100010100100110: color_data = 12'b111011101110;
20'b01001100010100100111: color_data = 12'b111011101110;
20'b01001100010100101000: color_data = 12'b111011101110;
20'b01001100010100101001: color_data = 12'b111011101110;
20'b01001100010100101010: color_data = 12'b111011101110;
20'b01001100010100101011: color_data = 12'b111011101110;
20'b01001100010100101100: color_data = 12'b111011101110;
20'b01001100010100101101: color_data = 12'b111011101110;
20'b01001100010100101111: color_data = 12'b111011101110;
20'b01001100010100110000: color_data = 12'b111011101110;
20'b01001100010100110001: color_data = 12'b111011101110;
20'b01001100010100110010: color_data = 12'b111011101110;
20'b01001100010100110011: color_data = 12'b111011101110;
20'b01001100010100110100: color_data = 12'b111011101110;
20'b01001100010100110101: color_data = 12'b111011101110;
20'b01001100010100110110: color_data = 12'b111011101110;
20'b01001100010100110111: color_data = 12'b111011101110;
20'b01001100010100111000: color_data = 12'b111011101110;
20'b01001100010101000100: color_data = 12'b111011101110;
20'b01001100010101000101: color_data = 12'b111011101110;
20'b01001100010101000110: color_data = 12'b111011101110;
20'b01001100010101000111: color_data = 12'b111011101110;
20'b01001100010101001000: color_data = 12'b111011101110;
20'b01001100010101001001: color_data = 12'b111011101110;
20'b01001100010101001010: color_data = 12'b111011101110;
20'b01001100010101001011: color_data = 12'b111011101110;
20'b01001100010101001100: color_data = 12'b111011101110;
20'b01001100010101001101: color_data = 12'b111011101110;
20'b01001100010101001111: color_data = 12'b111011101110;
20'b01001100010101010000: color_data = 12'b111011101110;
20'b01001100010101010001: color_data = 12'b111011101110;
20'b01001100010101010010: color_data = 12'b111011101110;
20'b01001100010101010011: color_data = 12'b111011101110;
20'b01001100010101010100: color_data = 12'b111011101110;
20'b01001100010101010101: color_data = 12'b111011101110;
20'b01001100010101010110: color_data = 12'b111011101110;
20'b01001100010101010111: color_data = 12'b111011101110;
20'b01001100010101011000: color_data = 12'b111011101110;
20'b01001100010110011100: color_data = 12'b111011101110;
20'b01001100010110011101: color_data = 12'b111011101110;
20'b01001100010110011110: color_data = 12'b111011101110;
20'b01001100010110011111: color_data = 12'b111011101110;
20'b01001100010110100000: color_data = 12'b111011101110;
20'b01001100010110100001: color_data = 12'b111011101110;
20'b01001100010110100010: color_data = 12'b111011101110;
20'b01001100010110100011: color_data = 12'b111011101110;
20'b01001100010110100100: color_data = 12'b111011101110;
20'b01001100010110100101: color_data = 12'b111011101110;
20'b01001100010110100111: color_data = 12'b111011101110;
20'b01001100010110101000: color_data = 12'b111011101110;
20'b01001100010110101001: color_data = 12'b111011101110;
20'b01001100010110101010: color_data = 12'b111011101110;
20'b01001100010110101011: color_data = 12'b111011101110;
20'b01001100010110101100: color_data = 12'b111011101110;
20'b01001100010110101101: color_data = 12'b111011101110;
20'b01001100010110101110: color_data = 12'b111011101110;
20'b01001100010110101111: color_data = 12'b111011101110;
20'b01001100010110110000: color_data = 12'b111011101110;
20'b01001100010110110010: color_data = 12'b111011101110;
20'b01001100010110110011: color_data = 12'b111011101110;
20'b01001100010110110100: color_data = 12'b111011101110;
20'b01001100010110110101: color_data = 12'b111011101110;
20'b01001100010110110110: color_data = 12'b111011101110;
20'b01001100010110110111: color_data = 12'b111011101110;
20'b01001100010110111000: color_data = 12'b111011101110;
20'b01001100010110111001: color_data = 12'b111011101110;
20'b01001100010110111010: color_data = 12'b111011101110;
20'b01001100010110111011: color_data = 12'b111011101110;
20'b01001100010110111101: color_data = 12'b111011101110;
20'b01001100010110111110: color_data = 12'b111011101110;
20'b01001100010110111111: color_data = 12'b111011101110;
20'b01001100010111000000: color_data = 12'b111011101110;
20'b01001100010111000001: color_data = 12'b111011101110;
20'b01001100010111000010: color_data = 12'b111011101110;
20'b01001100010111000011: color_data = 12'b111011101110;
20'b01001100010111000100: color_data = 12'b111011101110;
20'b01001100010111000101: color_data = 12'b111011101110;
20'b01001100010111000110: color_data = 12'b111011101110;
20'b01001100100010010110: color_data = 12'b111011101110;
20'b01001100100010010111: color_data = 12'b111011101110;
20'b01001100100010011000: color_data = 12'b111011101110;
20'b01001100100010011001: color_data = 12'b111011101110;
20'b01001100100010011010: color_data = 12'b111011101110;
20'b01001100100010011011: color_data = 12'b111011101110;
20'b01001100100010011100: color_data = 12'b111011101110;
20'b01001100100010011101: color_data = 12'b111011101110;
20'b01001100100010011110: color_data = 12'b111011101110;
20'b01001100100010011111: color_data = 12'b111011101110;
20'b01001100100010100001: color_data = 12'b111011101110;
20'b01001100100010100010: color_data = 12'b111011101110;
20'b01001100100010100011: color_data = 12'b111011101110;
20'b01001100100010100100: color_data = 12'b111011101110;
20'b01001100100010100101: color_data = 12'b111011101110;
20'b01001100100010100110: color_data = 12'b111011101110;
20'b01001100100010100111: color_data = 12'b111011101110;
20'b01001100100010101000: color_data = 12'b111011101110;
20'b01001100100010101001: color_data = 12'b111011101110;
20'b01001100100010101010: color_data = 12'b111011101110;
20'b01001100100011001101: color_data = 12'b111011101110;
20'b01001100100011001110: color_data = 12'b111011101110;
20'b01001100100011001111: color_data = 12'b111011101110;
20'b01001100100011010000: color_data = 12'b111011101110;
20'b01001100100011010001: color_data = 12'b111011101110;
20'b01001100100011010010: color_data = 12'b111011101110;
20'b01001100100011010011: color_data = 12'b111011101110;
20'b01001100100011010100: color_data = 12'b111011101110;
20'b01001100100011010101: color_data = 12'b111011101110;
20'b01001100100011010110: color_data = 12'b111011101110;
20'b01001100100011011000: color_data = 12'b111011101110;
20'b01001100100011011001: color_data = 12'b111011101110;
20'b01001100100011011010: color_data = 12'b111011101110;
20'b01001100100011011011: color_data = 12'b111011101110;
20'b01001100100011011100: color_data = 12'b111011101110;
20'b01001100100011011101: color_data = 12'b111011101110;
20'b01001100100011011110: color_data = 12'b111011101110;
20'b01001100100011011111: color_data = 12'b111011101110;
20'b01001100100011100000: color_data = 12'b111011101110;
20'b01001100100011100001: color_data = 12'b111011101110;
20'b01001100100011101101: color_data = 12'b111011101110;
20'b01001100100011101110: color_data = 12'b111011101110;
20'b01001100100011101111: color_data = 12'b111011101110;
20'b01001100100011110000: color_data = 12'b111011101110;
20'b01001100100011110001: color_data = 12'b111011101110;
20'b01001100100011110010: color_data = 12'b111011101110;
20'b01001100100011110011: color_data = 12'b111011101110;
20'b01001100100011110100: color_data = 12'b111011101110;
20'b01001100100011110101: color_data = 12'b111011101110;
20'b01001100100011110110: color_data = 12'b111011101110;
20'b01001100100011111000: color_data = 12'b111011101110;
20'b01001100100011111001: color_data = 12'b111011101110;
20'b01001100100011111010: color_data = 12'b111011101110;
20'b01001100100011111011: color_data = 12'b111011101110;
20'b01001100100011111100: color_data = 12'b111011101110;
20'b01001100100011111101: color_data = 12'b111011101110;
20'b01001100100011111110: color_data = 12'b111011101110;
20'b01001100100011111111: color_data = 12'b111011101110;
20'b01001100100100000000: color_data = 12'b111011101110;
20'b01001100100100000001: color_data = 12'b111011101110;
20'b01001100100100100100: color_data = 12'b111011101110;
20'b01001100100100100101: color_data = 12'b111011101110;
20'b01001100100100100110: color_data = 12'b111011101110;
20'b01001100100100100111: color_data = 12'b111011101110;
20'b01001100100100101000: color_data = 12'b111011101110;
20'b01001100100100101001: color_data = 12'b111011101110;
20'b01001100100100101010: color_data = 12'b111011101110;
20'b01001100100100101011: color_data = 12'b111011101110;
20'b01001100100100101100: color_data = 12'b111011101110;
20'b01001100100100101101: color_data = 12'b111011101110;
20'b01001100100100101111: color_data = 12'b111011101110;
20'b01001100100100110000: color_data = 12'b111011101110;
20'b01001100100100110001: color_data = 12'b111011101110;
20'b01001100100100110010: color_data = 12'b111011101110;
20'b01001100100100110011: color_data = 12'b111011101110;
20'b01001100100100110100: color_data = 12'b111011101110;
20'b01001100100100110101: color_data = 12'b111011101110;
20'b01001100100100110110: color_data = 12'b111011101110;
20'b01001100100100110111: color_data = 12'b111011101110;
20'b01001100100100111000: color_data = 12'b111011101110;
20'b01001100100101000100: color_data = 12'b111011101110;
20'b01001100100101000101: color_data = 12'b111011101110;
20'b01001100100101000110: color_data = 12'b111011101110;
20'b01001100100101000111: color_data = 12'b111011101110;
20'b01001100100101001000: color_data = 12'b111011101110;
20'b01001100100101001001: color_data = 12'b111011101110;
20'b01001100100101001010: color_data = 12'b111011101110;
20'b01001100100101001011: color_data = 12'b111011101110;
20'b01001100100101001100: color_data = 12'b111011101110;
20'b01001100100101001101: color_data = 12'b111011101110;
20'b01001100100101001111: color_data = 12'b111011101110;
20'b01001100100101010000: color_data = 12'b111011101110;
20'b01001100100101010001: color_data = 12'b111011101110;
20'b01001100100101010010: color_data = 12'b111011101110;
20'b01001100100101010011: color_data = 12'b111011101110;
20'b01001100100101010100: color_data = 12'b111011101110;
20'b01001100100101010101: color_data = 12'b111011101110;
20'b01001100100101010110: color_data = 12'b111011101110;
20'b01001100100101010111: color_data = 12'b111011101110;
20'b01001100100101011000: color_data = 12'b111011101110;
20'b01001100100110011100: color_data = 12'b111011101110;
20'b01001100100110011101: color_data = 12'b111011101110;
20'b01001100100110011110: color_data = 12'b111011101110;
20'b01001100100110011111: color_data = 12'b111011101110;
20'b01001100100110100000: color_data = 12'b111011101110;
20'b01001100100110100001: color_data = 12'b111011101110;
20'b01001100100110100010: color_data = 12'b111011101110;
20'b01001100100110100011: color_data = 12'b111011101110;
20'b01001100100110100100: color_data = 12'b111011101110;
20'b01001100100110100101: color_data = 12'b111011101110;
20'b01001100100110100111: color_data = 12'b111011101110;
20'b01001100100110101000: color_data = 12'b111011101110;
20'b01001100100110101001: color_data = 12'b111011101110;
20'b01001100100110101010: color_data = 12'b111011101110;
20'b01001100100110101011: color_data = 12'b111011101110;
20'b01001100100110101100: color_data = 12'b111011101110;
20'b01001100100110101101: color_data = 12'b111011101110;
20'b01001100100110101110: color_data = 12'b111011101110;
20'b01001100100110101111: color_data = 12'b111011101110;
20'b01001100100110110000: color_data = 12'b111011101110;
20'b01001100100110110010: color_data = 12'b111011101110;
20'b01001100100110110011: color_data = 12'b111011101110;
20'b01001100100110110100: color_data = 12'b111011101110;
20'b01001100100110110101: color_data = 12'b111011101110;
20'b01001100100110110110: color_data = 12'b111011101110;
20'b01001100100110110111: color_data = 12'b111011101110;
20'b01001100100110111000: color_data = 12'b111011101110;
20'b01001100100110111001: color_data = 12'b111011101110;
20'b01001100100110111010: color_data = 12'b111011101110;
20'b01001100100110111011: color_data = 12'b111011101110;
20'b01001100100110111101: color_data = 12'b111011101110;
20'b01001100100110111110: color_data = 12'b111011101110;
20'b01001100100110111111: color_data = 12'b111011101110;
20'b01001100100111000000: color_data = 12'b111011101110;
20'b01001100100111000001: color_data = 12'b111011101110;
20'b01001100100111000010: color_data = 12'b111011101110;
20'b01001100100111000011: color_data = 12'b111011101110;
20'b01001100100111000100: color_data = 12'b111011101110;
20'b01001100100111000101: color_data = 12'b111011101110;
20'b01001100100111000110: color_data = 12'b111011101110;
20'b01001100110010010110: color_data = 12'b111011101110;
20'b01001100110010010111: color_data = 12'b111011101110;
20'b01001100110010011000: color_data = 12'b111011101110;
20'b01001100110010011001: color_data = 12'b111011101110;
20'b01001100110010011010: color_data = 12'b111011101110;
20'b01001100110010011011: color_data = 12'b111011101110;
20'b01001100110010011100: color_data = 12'b111011101110;
20'b01001100110010011101: color_data = 12'b111011101110;
20'b01001100110010011110: color_data = 12'b111011101110;
20'b01001100110010011111: color_data = 12'b111011101110;
20'b01001100110010100001: color_data = 12'b111011101110;
20'b01001100110010100010: color_data = 12'b111011101110;
20'b01001100110010100011: color_data = 12'b111011101110;
20'b01001100110010100100: color_data = 12'b111011101110;
20'b01001100110010100101: color_data = 12'b111011101110;
20'b01001100110010100110: color_data = 12'b111011101110;
20'b01001100110010100111: color_data = 12'b111011101110;
20'b01001100110010101000: color_data = 12'b111011101110;
20'b01001100110010101001: color_data = 12'b111011101110;
20'b01001100110010101010: color_data = 12'b111011101110;
20'b01001100110011001101: color_data = 12'b111011101110;
20'b01001100110011001110: color_data = 12'b111011101110;
20'b01001100110011001111: color_data = 12'b111011101110;
20'b01001100110011010000: color_data = 12'b111011101110;
20'b01001100110011010001: color_data = 12'b111011101110;
20'b01001100110011010010: color_data = 12'b111011101110;
20'b01001100110011010011: color_data = 12'b111011101110;
20'b01001100110011010100: color_data = 12'b111011101110;
20'b01001100110011010101: color_data = 12'b111011101110;
20'b01001100110011010110: color_data = 12'b111011101110;
20'b01001100110011011000: color_data = 12'b111011101110;
20'b01001100110011011001: color_data = 12'b111011101110;
20'b01001100110011011010: color_data = 12'b111011101110;
20'b01001100110011011011: color_data = 12'b111011101110;
20'b01001100110011011100: color_data = 12'b111011101110;
20'b01001100110011011101: color_data = 12'b111011101110;
20'b01001100110011011110: color_data = 12'b111011101110;
20'b01001100110011011111: color_data = 12'b111011101110;
20'b01001100110011100000: color_data = 12'b111011101110;
20'b01001100110011100001: color_data = 12'b111011101110;
20'b01001100110011101101: color_data = 12'b111011101110;
20'b01001100110011101110: color_data = 12'b111011101110;
20'b01001100110011101111: color_data = 12'b111011101110;
20'b01001100110011110000: color_data = 12'b111011101110;
20'b01001100110011110001: color_data = 12'b111011101110;
20'b01001100110011110010: color_data = 12'b111011101110;
20'b01001100110011110011: color_data = 12'b111011101110;
20'b01001100110011110100: color_data = 12'b111011101110;
20'b01001100110011110101: color_data = 12'b111011101110;
20'b01001100110011110110: color_data = 12'b111011101110;
20'b01001100110011111000: color_data = 12'b111011101110;
20'b01001100110011111001: color_data = 12'b111011101110;
20'b01001100110011111010: color_data = 12'b111011101110;
20'b01001100110011111011: color_data = 12'b111011101110;
20'b01001100110011111100: color_data = 12'b111011101110;
20'b01001100110011111101: color_data = 12'b111011101110;
20'b01001100110011111110: color_data = 12'b111011101110;
20'b01001100110011111111: color_data = 12'b111011101110;
20'b01001100110100000000: color_data = 12'b111011101110;
20'b01001100110100000001: color_data = 12'b111011101110;
20'b01001100110100100100: color_data = 12'b111011101110;
20'b01001100110100100101: color_data = 12'b111011101110;
20'b01001100110100100110: color_data = 12'b111011101110;
20'b01001100110100100111: color_data = 12'b111011101110;
20'b01001100110100101000: color_data = 12'b111011101110;
20'b01001100110100101001: color_data = 12'b111011101110;
20'b01001100110100101010: color_data = 12'b111011101110;
20'b01001100110100101011: color_data = 12'b111011101110;
20'b01001100110100101100: color_data = 12'b111011101110;
20'b01001100110100101101: color_data = 12'b111011101110;
20'b01001100110100101111: color_data = 12'b111011101110;
20'b01001100110100110000: color_data = 12'b111011101110;
20'b01001100110100110001: color_data = 12'b111011101110;
20'b01001100110100110010: color_data = 12'b111011101110;
20'b01001100110100110011: color_data = 12'b111011101110;
20'b01001100110100110100: color_data = 12'b111011101110;
20'b01001100110100110101: color_data = 12'b111011101110;
20'b01001100110100110110: color_data = 12'b111011101110;
20'b01001100110100110111: color_data = 12'b111011101110;
20'b01001100110100111000: color_data = 12'b111011101110;
20'b01001100110101000100: color_data = 12'b111011101110;
20'b01001100110101000101: color_data = 12'b111011101110;
20'b01001100110101000110: color_data = 12'b111011101110;
20'b01001100110101000111: color_data = 12'b111011101110;
20'b01001100110101001000: color_data = 12'b111011101110;
20'b01001100110101001001: color_data = 12'b111011101110;
20'b01001100110101001010: color_data = 12'b111011101110;
20'b01001100110101001011: color_data = 12'b111011101110;
20'b01001100110101001100: color_data = 12'b111011101110;
20'b01001100110101001101: color_data = 12'b111011101110;
20'b01001100110101001111: color_data = 12'b111011101110;
20'b01001100110101010000: color_data = 12'b111011101110;
20'b01001100110101010001: color_data = 12'b111011101110;
20'b01001100110101010010: color_data = 12'b111011101110;
20'b01001100110101010011: color_data = 12'b111011101110;
20'b01001100110101010100: color_data = 12'b111011101110;
20'b01001100110101010101: color_data = 12'b111011101110;
20'b01001100110101010110: color_data = 12'b111011101110;
20'b01001100110101010111: color_data = 12'b111011101110;
20'b01001100110101011000: color_data = 12'b111011101110;
20'b01001100110110011100: color_data = 12'b111011101110;
20'b01001100110110011101: color_data = 12'b111011101110;
20'b01001100110110011110: color_data = 12'b111011101110;
20'b01001100110110011111: color_data = 12'b111011101110;
20'b01001100110110100000: color_data = 12'b111011101110;
20'b01001100110110100001: color_data = 12'b111011101110;
20'b01001100110110100010: color_data = 12'b111011101110;
20'b01001100110110100011: color_data = 12'b111011101110;
20'b01001100110110100100: color_data = 12'b111011101110;
20'b01001100110110100101: color_data = 12'b111011101110;
20'b01001100110110100111: color_data = 12'b111011101110;
20'b01001100110110101000: color_data = 12'b111011101110;
20'b01001100110110101001: color_data = 12'b111011101110;
20'b01001100110110101010: color_data = 12'b111011101110;
20'b01001100110110101011: color_data = 12'b111011101110;
20'b01001100110110101100: color_data = 12'b111011101110;
20'b01001100110110101101: color_data = 12'b111011101110;
20'b01001100110110101110: color_data = 12'b111011101110;
20'b01001100110110101111: color_data = 12'b111011101110;
20'b01001100110110110000: color_data = 12'b111011101110;
20'b01001100110110110010: color_data = 12'b111011101110;
20'b01001100110110110011: color_data = 12'b111011101110;
20'b01001100110110110100: color_data = 12'b111011101110;
20'b01001100110110110101: color_data = 12'b111011101110;
20'b01001100110110110110: color_data = 12'b111011101110;
20'b01001100110110110111: color_data = 12'b111011101110;
20'b01001100110110111000: color_data = 12'b111011101110;
20'b01001100110110111001: color_data = 12'b111011101110;
20'b01001100110110111010: color_data = 12'b111011101110;
20'b01001100110110111011: color_data = 12'b111011101110;
20'b01001100110110111101: color_data = 12'b111011101110;
20'b01001100110110111110: color_data = 12'b111011101110;
20'b01001100110110111111: color_data = 12'b111011101110;
20'b01001100110111000000: color_data = 12'b111011101110;
20'b01001100110111000001: color_data = 12'b111011101110;
20'b01001100110111000010: color_data = 12'b111011101110;
20'b01001100110111000011: color_data = 12'b111011101110;
20'b01001100110111000100: color_data = 12'b111011101110;
20'b01001100110111000101: color_data = 12'b111011101110;
20'b01001100110111000110: color_data = 12'b111011101110;
20'b01001101000010010110: color_data = 12'b111011101110;
20'b01001101000010010111: color_data = 12'b111011101110;
20'b01001101000010011000: color_data = 12'b111011101110;
20'b01001101000010011001: color_data = 12'b111011101110;
20'b01001101000010011010: color_data = 12'b111011101110;
20'b01001101000010011011: color_data = 12'b111011101110;
20'b01001101000010011100: color_data = 12'b111011101110;
20'b01001101000010011101: color_data = 12'b111011101110;
20'b01001101000010011110: color_data = 12'b111011101110;
20'b01001101000010011111: color_data = 12'b111011101110;
20'b01001101000010100001: color_data = 12'b111011101110;
20'b01001101000010100010: color_data = 12'b111011101110;
20'b01001101000010100011: color_data = 12'b111011101110;
20'b01001101000010100100: color_data = 12'b111011101110;
20'b01001101000010100101: color_data = 12'b111011101110;
20'b01001101000010100110: color_data = 12'b111011101110;
20'b01001101000010100111: color_data = 12'b111011101110;
20'b01001101000010101000: color_data = 12'b111011101110;
20'b01001101000010101001: color_data = 12'b111011101110;
20'b01001101000010101010: color_data = 12'b111011101110;
20'b01001101000011001101: color_data = 12'b111011101110;
20'b01001101000011001110: color_data = 12'b111011101110;
20'b01001101000011001111: color_data = 12'b111011101110;
20'b01001101000011010000: color_data = 12'b111011101110;
20'b01001101000011010001: color_data = 12'b111011101110;
20'b01001101000011010010: color_data = 12'b111011101110;
20'b01001101000011010011: color_data = 12'b111011101110;
20'b01001101000011010100: color_data = 12'b111011101110;
20'b01001101000011010101: color_data = 12'b111011101110;
20'b01001101000011010110: color_data = 12'b111011101110;
20'b01001101000011011000: color_data = 12'b111011101110;
20'b01001101000011011001: color_data = 12'b111011101110;
20'b01001101000011011010: color_data = 12'b111011101110;
20'b01001101000011011011: color_data = 12'b111011101110;
20'b01001101000011011100: color_data = 12'b111011101110;
20'b01001101000011011101: color_data = 12'b111011101110;
20'b01001101000011011110: color_data = 12'b111011101110;
20'b01001101000011011111: color_data = 12'b111011101110;
20'b01001101000011100000: color_data = 12'b111011101110;
20'b01001101000011100001: color_data = 12'b111011101110;
20'b01001101000011101101: color_data = 12'b111011101110;
20'b01001101000011101110: color_data = 12'b111011101110;
20'b01001101000011101111: color_data = 12'b111011101110;
20'b01001101000011110000: color_data = 12'b111011101110;
20'b01001101000011110001: color_data = 12'b111011101110;
20'b01001101000011110010: color_data = 12'b111011101110;
20'b01001101000011110011: color_data = 12'b111011101110;
20'b01001101000011110100: color_data = 12'b111011101110;
20'b01001101000011110101: color_data = 12'b111011101110;
20'b01001101000011110110: color_data = 12'b111011101110;
20'b01001101000011111000: color_data = 12'b111011101110;
20'b01001101000011111001: color_data = 12'b111011101110;
20'b01001101000011111010: color_data = 12'b111011101110;
20'b01001101000011111011: color_data = 12'b111011101110;
20'b01001101000011111100: color_data = 12'b111011101110;
20'b01001101000011111101: color_data = 12'b111011101110;
20'b01001101000011111110: color_data = 12'b111011101110;
20'b01001101000011111111: color_data = 12'b111011101110;
20'b01001101000100000000: color_data = 12'b111011101110;
20'b01001101000100000001: color_data = 12'b111011101110;
20'b01001101000100100100: color_data = 12'b111011101110;
20'b01001101000100100101: color_data = 12'b111011101110;
20'b01001101000100100110: color_data = 12'b111011101110;
20'b01001101000100100111: color_data = 12'b111011101110;
20'b01001101000100101000: color_data = 12'b111011101110;
20'b01001101000100101001: color_data = 12'b111011101110;
20'b01001101000100101010: color_data = 12'b111011101110;
20'b01001101000100101011: color_data = 12'b111011101110;
20'b01001101000100101100: color_data = 12'b111011101110;
20'b01001101000100101101: color_data = 12'b111011101110;
20'b01001101000100101111: color_data = 12'b111011101110;
20'b01001101000100110000: color_data = 12'b111011101110;
20'b01001101000100110001: color_data = 12'b111011101110;
20'b01001101000100110010: color_data = 12'b111011101110;
20'b01001101000100110011: color_data = 12'b111011101110;
20'b01001101000100110100: color_data = 12'b111011101110;
20'b01001101000100110101: color_data = 12'b111011101110;
20'b01001101000100110110: color_data = 12'b111011101110;
20'b01001101000100110111: color_data = 12'b111011101110;
20'b01001101000100111000: color_data = 12'b111011101110;
20'b01001101000101000100: color_data = 12'b111011101110;
20'b01001101000101000101: color_data = 12'b111011101110;
20'b01001101000101000110: color_data = 12'b111011101110;
20'b01001101000101000111: color_data = 12'b111011101110;
20'b01001101000101001000: color_data = 12'b111011101110;
20'b01001101000101001001: color_data = 12'b111011101110;
20'b01001101000101001010: color_data = 12'b111011101110;
20'b01001101000101001011: color_data = 12'b111011101110;
20'b01001101000101001100: color_data = 12'b111011101110;
20'b01001101000101001101: color_data = 12'b111011101110;
20'b01001101000101001111: color_data = 12'b111011101110;
20'b01001101000101010000: color_data = 12'b111011101110;
20'b01001101000101010001: color_data = 12'b111011101110;
20'b01001101000101010010: color_data = 12'b111011101110;
20'b01001101000101010011: color_data = 12'b111011101110;
20'b01001101000101010100: color_data = 12'b111011101110;
20'b01001101000101010101: color_data = 12'b111011101110;
20'b01001101000101010110: color_data = 12'b111011101110;
20'b01001101000101010111: color_data = 12'b111011101110;
20'b01001101000101011000: color_data = 12'b111011101110;
20'b01001101000110011100: color_data = 12'b111011101110;
20'b01001101000110011101: color_data = 12'b111011101110;
20'b01001101000110011110: color_data = 12'b111011101110;
20'b01001101000110011111: color_data = 12'b111011101110;
20'b01001101000110100000: color_data = 12'b111011101110;
20'b01001101000110100001: color_data = 12'b111011101110;
20'b01001101000110100010: color_data = 12'b111011101110;
20'b01001101000110100011: color_data = 12'b111011101110;
20'b01001101000110100100: color_data = 12'b111011101110;
20'b01001101000110100101: color_data = 12'b111011101110;
20'b01001101000110100111: color_data = 12'b111011101110;
20'b01001101000110101000: color_data = 12'b111011101110;
20'b01001101000110101001: color_data = 12'b111011101110;
20'b01001101000110101010: color_data = 12'b111011101110;
20'b01001101000110101011: color_data = 12'b111011101110;
20'b01001101000110101100: color_data = 12'b111011101110;
20'b01001101000110101101: color_data = 12'b111011101110;
20'b01001101000110101110: color_data = 12'b111011101110;
20'b01001101000110101111: color_data = 12'b111011101110;
20'b01001101000110110000: color_data = 12'b111011101110;
20'b01001101000110110010: color_data = 12'b111011101110;
20'b01001101000110110011: color_data = 12'b111011101110;
20'b01001101000110110100: color_data = 12'b111011101110;
20'b01001101000110110101: color_data = 12'b111011101110;
20'b01001101000110110110: color_data = 12'b111011101110;
20'b01001101000110110111: color_data = 12'b111011101110;
20'b01001101000110111000: color_data = 12'b111011101110;
20'b01001101000110111001: color_data = 12'b111011101110;
20'b01001101000110111010: color_data = 12'b111011101110;
20'b01001101000110111011: color_data = 12'b111011101110;
20'b01001101000110111101: color_data = 12'b111011101110;
20'b01001101000110111110: color_data = 12'b111011101110;
20'b01001101000110111111: color_data = 12'b111011101110;
20'b01001101000111000000: color_data = 12'b111011101110;
20'b01001101000111000001: color_data = 12'b111011101110;
20'b01001101000111000010: color_data = 12'b111011101110;
20'b01001101000111000011: color_data = 12'b111011101110;
20'b01001101000111000100: color_data = 12'b111011101110;
20'b01001101000111000101: color_data = 12'b111011101110;
20'b01001101000111000110: color_data = 12'b111011101110;
20'b01001101010010010110: color_data = 12'b111011101110;
20'b01001101010010010111: color_data = 12'b111011101110;
20'b01001101010010011000: color_data = 12'b111011101110;
20'b01001101010010011001: color_data = 12'b111011101110;
20'b01001101010010011010: color_data = 12'b111011101110;
20'b01001101010010011011: color_data = 12'b111011101110;
20'b01001101010010011100: color_data = 12'b111011101110;
20'b01001101010010011101: color_data = 12'b111011101110;
20'b01001101010010011110: color_data = 12'b111011101110;
20'b01001101010010011111: color_data = 12'b111011101110;
20'b01001101010010100001: color_data = 12'b111011101110;
20'b01001101010010100010: color_data = 12'b111011101110;
20'b01001101010010100011: color_data = 12'b111011101110;
20'b01001101010010100100: color_data = 12'b111011101110;
20'b01001101010010100101: color_data = 12'b111011101110;
20'b01001101010010100110: color_data = 12'b111011101110;
20'b01001101010010100111: color_data = 12'b111011101110;
20'b01001101010010101000: color_data = 12'b111011101110;
20'b01001101010010101001: color_data = 12'b111011101110;
20'b01001101010010101010: color_data = 12'b111011101110;
20'b01001101010011001101: color_data = 12'b111011101110;
20'b01001101010011001110: color_data = 12'b111011101110;
20'b01001101010011001111: color_data = 12'b111011101110;
20'b01001101010011010000: color_data = 12'b111011101110;
20'b01001101010011010001: color_data = 12'b111011101110;
20'b01001101010011010010: color_data = 12'b111011101110;
20'b01001101010011010011: color_data = 12'b111011101110;
20'b01001101010011010100: color_data = 12'b111011101110;
20'b01001101010011010101: color_data = 12'b111011101110;
20'b01001101010011010110: color_data = 12'b111011101110;
20'b01001101010011011000: color_data = 12'b111011101110;
20'b01001101010011011001: color_data = 12'b111011101110;
20'b01001101010011011010: color_data = 12'b111011101110;
20'b01001101010011011011: color_data = 12'b111011101110;
20'b01001101010011011100: color_data = 12'b111011101110;
20'b01001101010011011101: color_data = 12'b111011101110;
20'b01001101010011011110: color_data = 12'b111011101110;
20'b01001101010011011111: color_data = 12'b111011101110;
20'b01001101010011100000: color_data = 12'b111011101110;
20'b01001101010011100001: color_data = 12'b111011101110;
20'b01001101010011101101: color_data = 12'b111011101110;
20'b01001101010011101110: color_data = 12'b111011101110;
20'b01001101010011101111: color_data = 12'b111011101110;
20'b01001101010011110000: color_data = 12'b111011101110;
20'b01001101010011110001: color_data = 12'b111011101110;
20'b01001101010011110010: color_data = 12'b111011101110;
20'b01001101010011110011: color_data = 12'b111011101110;
20'b01001101010011110100: color_data = 12'b111011101110;
20'b01001101010011110101: color_data = 12'b111011101110;
20'b01001101010011110110: color_data = 12'b111011101110;
20'b01001101010011111000: color_data = 12'b111011101110;
20'b01001101010011111001: color_data = 12'b111011101110;
20'b01001101010011111010: color_data = 12'b111011101110;
20'b01001101010011111011: color_data = 12'b111011101110;
20'b01001101010011111100: color_data = 12'b111011101110;
20'b01001101010011111101: color_data = 12'b111011101110;
20'b01001101010011111110: color_data = 12'b111011101110;
20'b01001101010011111111: color_data = 12'b111011101110;
20'b01001101010100000000: color_data = 12'b111011101110;
20'b01001101010100000001: color_data = 12'b111011101110;
20'b01001101010100100100: color_data = 12'b111011101110;
20'b01001101010100100101: color_data = 12'b111011101110;
20'b01001101010100100110: color_data = 12'b111011101110;
20'b01001101010100100111: color_data = 12'b111011101110;
20'b01001101010100101000: color_data = 12'b111011101110;
20'b01001101010100101001: color_data = 12'b111011101110;
20'b01001101010100101010: color_data = 12'b111011101110;
20'b01001101010100101011: color_data = 12'b111011101110;
20'b01001101010100101100: color_data = 12'b111011101110;
20'b01001101010100101101: color_data = 12'b111011101110;
20'b01001101010100101111: color_data = 12'b111011101110;
20'b01001101010100110000: color_data = 12'b111011101110;
20'b01001101010100110001: color_data = 12'b111011101110;
20'b01001101010100110010: color_data = 12'b111011101110;
20'b01001101010100110011: color_data = 12'b111011101110;
20'b01001101010100110100: color_data = 12'b111011101110;
20'b01001101010100110101: color_data = 12'b111011101110;
20'b01001101010100110110: color_data = 12'b111011101110;
20'b01001101010100110111: color_data = 12'b111011101110;
20'b01001101010100111000: color_data = 12'b111011101110;
20'b01001101010101000100: color_data = 12'b111011101110;
20'b01001101010101000101: color_data = 12'b111011101110;
20'b01001101010101000110: color_data = 12'b111011101110;
20'b01001101010101000111: color_data = 12'b111011101110;
20'b01001101010101001000: color_data = 12'b111011101110;
20'b01001101010101001001: color_data = 12'b111011101110;
20'b01001101010101001010: color_data = 12'b111011101110;
20'b01001101010101001011: color_data = 12'b111011101110;
20'b01001101010101001100: color_data = 12'b111011101110;
20'b01001101010101001101: color_data = 12'b111011101110;
20'b01001101010101001111: color_data = 12'b111011101110;
20'b01001101010101010000: color_data = 12'b111011101110;
20'b01001101010101010001: color_data = 12'b111011101110;
20'b01001101010101010010: color_data = 12'b111011101110;
20'b01001101010101010011: color_data = 12'b111011101110;
20'b01001101010101010100: color_data = 12'b111011101110;
20'b01001101010101010101: color_data = 12'b111011101110;
20'b01001101010101010110: color_data = 12'b111011101110;
20'b01001101010101010111: color_data = 12'b111011101110;
20'b01001101010101011000: color_data = 12'b111011101110;
20'b01001101010110011100: color_data = 12'b111011101110;
20'b01001101010110011101: color_data = 12'b111011101110;
20'b01001101010110011110: color_data = 12'b111011101110;
20'b01001101010110011111: color_data = 12'b111011101110;
20'b01001101010110100000: color_data = 12'b111011101110;
20'b01001101010110100001: color_data = 12'b111011101110;
20'b01001101010110100010: color_data = 12'b111011101110;
20'b01001101010110100011: color_data = 12'b111011101110;
20'b01001101010110100100: color_data = 12'b111011101110;
20'b01001101010110100101: color_data = 12'b111011101110;
20'b01001101010110100111: color_data = 12'b111011101110;
20'b01001101010110101000: color_data = 12'b111011101110;
20'b01001101010110101001: color_data = 12'b111011101110;
20'b01001101010110101010: color_data = 12'b111011101110;
20'b01001101010110101011: color_data = 12'b111011101110;
20'b01001101010110101100: color_data = 12'b111011101110;
20'b01001101010110101101: color_data = 12'b111011101110;
20'b01001101010110101110: color_data = 12'b111011101110;
20'b01001101010110101111: color_data = 12'b111011101110;
20'b01001101010110110000: color_data = 12'b111011101110;
20'b01001101010110110010: color_data = 12'b111011101110;
20'b01001101010110110011: color_data = 12'b111011101110;
20'b01001101010110110100: color_data = 12'b111011101110;
20'b01001101010110110101: color_data = 12'b111011101110;
20'b01001101010110110110: color_data = 12'b111011101110;
20'b01001101010110110111: color_data = 12'b111011101110;
20'b01001101010110111000: color_data = 12'b111011101110;
20'b01001101010110111001: color_data = 12'b111011101110;
20'b01001101010110111010: color_data = 12'b111011101110;
20'b01001101010110111011: color_data = 12'b111011101110;
20'b01001101010110111101: color_data = 12'b111011101110;
20'b01001101010110111110: color_data = 12'b111011101110;
20'b01001101010110111111: color_data = 12'b111011101110;
20'b01001101010111000000: color_data = 12'b111011101110;
20'b01001101010111000001: color_data = 12'b111011101110;
20'b01001101010111000010: color_data = 12'b111011101110;
20'b01001101010111000011: color_data = 12'b111011101110;
20'b01001101010111000100: color_data = 12'b111011101110;
20'b01001101010111000101: color_data = 12'b111011101110;
20'b01001101010111000110: color_data = 12'b111011101110;
20'b01001101110010010110: color_data = 12'b111011101110;
20'b01001101110010010111: color_data = 12'b111011101110;
20'b01001101110010011000: color_data = 12'b111011101110;
20'b01001101110010011001: color_data = 12'b111011101110;
20'b01001101110010011010: color_data = 12'b111011101110;
20'b01001101110010011011: color_data = 12'b111011101110;
20'b01001101110010011100: color_data = 12'b111011101110;
20'b01001101110010011101: color_data = 12'b111011101110;
20'b01001101110010011110: color_data = 12'b111011101110;
20'b01001101110010011111: color_data = 12'b111011101110;
20'b01001101110010100001: color_data = 12'b111011101110;
20'b01001101110010100010: color_data = 12'b111011101110;
20'b01001101110010100011: color_data = 12'b111011101110;
20'b01001101110010100100: color_data = 12'b111011101110;
20'b01001101110010100101: color_data = 12'b111011101110;
20'b01001101110010100110: color_data = 12'b111011101110;
20'b01001101110010100111: color_data = 12'b111011101110;
20'b01001101110010101000: color_data = 12'b111011101110;
20'b01001101110010101001: color_data = 12'b111011101110;
20'b01001101110010101010: color_data = 12'b111011101110;
20'b01001101110011001101: color_data = 12'b111011101110;
20'b01001101110011001110: color_data = 12'b111011101110;
20'b01001101110011001111: color_data = 12'b111011101110;
20'b01001101110011010000: color_data = 12'b111011101110;
20'b01001101110011010001: color_data = 12'b111011101110;
20'b01001101110011010010: color_data = 12'b111011101110;
20'b01001101110011010011: color_data = 12'b111011101110;
20'b01001101110011010100: color_data = 12'b111011101110;
20'b01001101110011010101: color_data = 12'b111011101110;
20'b01001101110011010110: color_data = 12'b111011101110;
20'b01001101110011011000: color_data = 12'b111011101110;
20'b01001101110011011001: color_data = 12'b111011101110;
20'b01001101110011011010: color_data = 12'b111011101110;
20'b01001101110011011011: color_data = 12'b111011101110;
20'b01001101110011011100: color_data = 12'b111011101110;
20'b01001101110011011101: color_data = 12'b111011101110;
20'b01001101110011011110: color_data = 12'b111011101110;
20'b01001101110011011111: color_data = 12'b111011101110;
20'b01001101110011100000: color_data = 12'b111011101110;
20'b01001101110011100001: color_data = 12'b111011101110;
20'b01001101110011101101: color_data = 12'b111011101110;
20'b01001101110011101110: color_data = 12'b111011101110;
20'b01001101110011101111: color_data = 12'b111011101110;
20'b01001101110011110000: color_data = 12'b111011101110;
20'b01001101110011110001: color_data = 12'b111011101110;
20'b01001101110011110010: color_data = 12'b111011101110;
20'b01001101110011110011: color_data = 12'b111011101110;
20'b01001101110011110100: color_data = 12'b111011101110;
20'b01001101110011110101: color_data = 12'b111011101110;
20'b01001101110011110110: color_data = 12'b111011101110;
20'b01001101110011111000: color_data = 12'b111011101110;
20'b01001101110011111001: color_data = 12'b111011101110;
20'b01001101110011111010: color_data = 12'b111011101110;
20'b01001101110011111011: color_data = 12'b111011101110;
20'b01001101110011111100: color_data = 12'b111011101110;
20'b01001101110011111101: color_data = 12'b111011101110;
20'b01001101110011111110: color_data = 12'b111011101110;
20'b01001101110011111111: color_data = 12'b111011101110;
20'b01001101110100000000: color_data = 12'b111011101110;
20'b01001101110100000001: color_data = 12'b111011101110;
20'b01001101110100000011: color_data = 12'b111011101110;
20'b01001101110100000100: color_data = 12'b111011101110;
20'b01001101110100000101: color_data = 12'b111011101110;
20'b01001101110100000110: color_data = 12'b111011101110;
20'b01001101110100000111: color_data = 12'b111011101110;
20'b01001101110100001000: color_data = 12'b111011101110;
20'b01001101110100001001: color_data = 12'b111011101110;
20'b01001101110100001010: color_data = 12'b111011101110;
20'b01001101110100001011: color_data = 12'b111011101110;
20'b01001101110100001100: color_data = 12'b111011101110;
20'b01001101110100011001: color_data = 12'b111011101110;
20'b01001101110100011010: color_data = 12'b111011101110;
20'b01001101110100011011: color_data = 12'b111011101110;
20'b01001101110100011100: color_data = 12'b111011101110;
20'b01001101110100011101: color_data = 12'b111011101110;
20'b01001101110100011110: color_data = 12'b111011101110;
20'b01001101110100011111: color_data = 12'b111011101110;
20'b01001101110100100000: color_data = 12'b111011101110;
20'b01001101110100100001: color_data = 12'b111011101110;
20'b01001101110100100010: color_data = 12'b111011101110;
20'b01001101110100100100: color_data = 12'b111011101110;
20'b01001101110100100101: color_data = 12'b111011101110;
20'b01001101110100100110: color_data = 12'b111011101110;
20'b01001101110100100111: color_data = 12'b111011101110;
20'b01001101110100101000: color_data = 12'b111011101110;
20'b01001101110100101001: color_data = 12'b111011101110;
20'b01001101110100101010: color_data = 12'b111011101110;
20'b01001101110100101011: color_data = 12'b111011101110;
20'b01001101110100101100: color_data = 12'b111011101110;
20'b01001101110100101101: color_data = 12'b111011101110;
20'b01001101110100101111: color_data = 12'b111011101110;
20'b01001101110100110000: color_data = 12'b111011101110;
20'b01001101110100110001: color_data = 12'b111011101110;
20'b01001101110100110010: color_data = 12'b111011101110;
20'b01001101110100110011: color_data = 12'b111011101110;
20'b01001101110100110100: color_data = 12'b111011101110;
20'b01001101110100110101: color_data = 12'b111011101110;
20'b01001101110100110110: color_data = 12'b111011101110;
20'b01001101110100110111: color_data = 12'b111011101110;
20'b01001101110100111000: color_data = 12'b111011101110;
20'b01001101110101000100: color_data = 12'b111011101110;
20'b01001101110101000101: color_data = 12'b111011101110;
20'b01001101110101000110: color_data = 12'b111011101110;
20'b01001101110101000111: color_data = 12'b111011101110;
20'b01001101110101001000: color_data = 12'b111011101110;
20'b01001101110101001001: color_data = 12'b111011101110;
20'b01001101110101001010: color_data = 12'b111011101110;
20'b01001101110101001011: color_data = 12'b111011101110;
20'b01001101110101001100: color_data = 12'b111011101110;
20'b01001101110101001101: color_data = 12'b111011101110;
20'b01001101110101001111: color_data = 12'b111011101110;
20'b01001101110101010000: color_data = 12'b111011101110;
20'b01001101110101010001: color_data = 12'b111011101110;
20'b01001101110101010010: color_data = 12'b111011101110;
20'b01001101110101010011: color_data = 12'b111011101110;
20'b01001101110101010100: color_data = 12'b111011101110;
20'b01001101110101010101: color_data = 12'b111011101110;
20'b01001101110101010110: color_data = 12'b111011101110;
20'b01001101110101010111: color_data = 12'b111011101110;
20'b01001101110101011000: color_data = 12'b111011101110;
20'b01001101110110011100: color_data = 12'b111011101110;
20'b01001101110110011101: color_data = 12'b111011101110;
20'b01001101110110011110: color_data = 12'b111011101110;
20'b01001101110110011111: color_data = 12'b111011101110;
20'b01001101110110100000: color_data = 12'b111011101110;
20'b01001101110110100001: color_data = 12'b111011101110;
20'b01001101110110100010: color_data = 12'b111011101110;
20'b01001101110110100011: color_data = 12'b111011101110;
20'b01001101110110100100: color_data = 12'b111011101110;
20'b01001101110110100101: color_data = 12'b111011101110;
20'b01001101110110100111: color_data = 12'b111011101110;
20'b01001101110110101000: color_data = 12'b111011101110;
20'b01001101110110101001: color_data = 12'b111011101110;
20'b01001101110110101010: color_data = 12'b111011101110;
20'b01001101110110101011: color_data = 12'b111011101110;
20'b01001101110110101100: color_data = 12'b111011101110;
20'b01001101110110101101: color_data = 12'b111011101110;
20'b01001101110110101110: color_data = 12'b111011101110;
20'b01001101110110101111: color_data = 12'b111011101110;
20'b01001101110110110000: color_data = 12'b111011101110;
20'b01001101110110111101: color_data = 12'b111011101110;
20'b01001101110110111110: color_data = 12'b111011101110;
20'b01001101110110111111: color_data = 12'b111011101110;
20'b01001101110111000000: color_data = 12'b111011101110;
20'b01001101110111000001: color_data = 12'b111011101110;
20'b01001101110111000010: color_data = 12'b111011101110;
20'b01001101110111000011: color_data = 12'b111011101110;
20'b01001101110111000100: color_data = 12'b111011101110;
20'b01001101110111000101: color_data = 12'b111011101110;
20'b01001101110111000110: color_data = 12'b111011101110;
20'b01001101110111001000: color_data = 12'b111011101110;
20'b01001101110111001001: color_data = 12'b111011101110;
20'b01001101110111001010: color_data = 12'b111011101110;
20'b01001101110111001011: color_data = 12'b111011101110;
20'b01001101110111001100: color_data = 12'b111011101110;
20'b01001101110111001101: color_data = 12'b111011101110;
20'b01001101110111001110: color_data = 12'b111011101110;
20'b01001101110111001111: color_data = 12'b111011101110;
20'b01001101110111010000: color_data = 12'b111011101110;
20'b01001101110111010001: color_data = 12'b111011101110;
20'b01001110000010010110: color_data = 12'b111011101110;
20'b01001110000010010111: color_data = 12'b111011101110;
20'b01001110000010011000: color_data = 12'b111011101110;
20'b01001110000010011001: color_data = 12'b111011101110;
20'b01001110000010011010: color_data = 12'b111011101110;
20'b01001110000010011011: color_data = 12'b111011101110;
20'b01001110000010011100: color_data = 12'b111011101110;
20'b01001110000010011101: color_data = 12'b111011101110;
20'b01001110000010011110: color_data = 12'b111011101110;
20'b01001110000010011111: color_data = 12'b111011101110;
20'b01001110000010100001: color_data = 12'b111011101110;
20'b01001110000010100010: color_data = 12'b111011101110;
20'b01001110000010100011: color_data = 12'b111011101110;
20'b01001110000010100100: color_data = 12'b111011101110;
20'b01001110000010100101: color_data = 12'b111011101110;
20'b01001110000010100110: color_data = 12'b111011101110;
20'b01001110000010100111: color_data = 12'b111011101110;
20'b01001110000010101000: color_data = 12'b111011101110;
20'b01001110000010101001: color_data = 12'b111011101110;
20'b01001110000010101010: color_data = 12'b111011101110;
20'b01001110000011001101: color_data = 12'b111011101110;
20'b01001110000011001110: color_data = 12'b111011101110;
20'b01001110000011001111: color_data = 12'b111011101110;
20'b01001110000011010000: color_data = 12'b111011101110;
20'b01001110000011010001: color_data = 12'b111011101110;
20'b01001110000011010010: color_data = 12'b111011101110;
20'b01001110000011010011: color_data = 12'b111011101110;
20'b01001110000011010100: color_data = 12'b111011101110;
20'b01001110000011010101: color_data = 12'b111011101110;
20'b01001110000011010110: color_data = 12'b111011101110;
20'b01001110000011011000: color_data = 12'b111011101110;
20'b01001110000011011001: color_data = 12'b111011101110;
20'b01001110000011011010: color_data = 12'b111011101110;
20'b01001110000011011011: color_data = 12'b111011101110;
20'b01001110000011011100: color_data = 12'b111011101110;
20'b01001110000011011101: color_data = 12'b111011101110;
20'b01001110000011011110: color_data = 12'b111011101110;
20'b01001110000011011111: color_data = 12'b111011101110;
20'b01001110000011100000: color_data = 12'b111011101110;
20'b01001110000011100001: color_data = 12'b111011101110;
20'b01001110000011101101: color_data = 12'b111011101110;
20'b01001110000011101110: color_data = 12'b111011101110;
20'b01001110000011101111: color_data = 12'b111011101110;
20'b01001110000011110000: color_data = 12'b111011101110;
20'b01001110000011110001: color_data = 12'b111011101110;
20'b01001110000011110010: color_data = 12'b111011101110;
20'b01001110000011110011: color_data = 12'b111011101110;
20'b01001110000011110100: color_data = 12'b111011101110;
20'b01001110000011110101: color_data = 12'b111011101110;
20'b01001110000011110110: color_data = 12'b111011101110;
20'b01001110000011111000: color_data = 12'b111011101110;
20'b01001110000011111001: color_data = 12'b111011101110;
20'b01001110000011111010: color_data = 12'b111011101110;
20'b01001110000011111011: color_data = 12'b111011101110;
20'b01001110000011111100: color_data = 12'b111011101110;
20'b01001110000011111101: color_data = 12'b111011101110;
20'b01001110000011111110: color_data = 12'b111011101110;
20'b01001110000011111111: color_data = 12'b111011101110;
20'b01001110000100000000: color_data = 12'b111011101110;
20'b01001110000100000001: color_data = 12'b111011101110;
20'b01001110000100000011: color_data = 12'b111011101110;
20'b01001110000100000100: color_data = 12'b111011101110;
20'b01001110000100000101: color_data = 12'b111011101110;
20'b01001110000100000110: color_data = 12'b111011101110;
20'b01001110000100000111: color_data = 12'b111011101110;
20'b01001110000100001000: color_data = 12'b111011101110;
20'b01001110000100001001: color_data = 12'b111011101110;
20'b01001110000100001010: color_data = 12'b111011101110;
20'b01001110000100001011: color_data = 12'b111011101110;
20'b01001110000100001100: color_data = 12'b111011101110;
20'b01001110000100011001: color_data = 12'b111011101110;
20'b01001110000100011010: color_data = 12'b111011101110;
20'b01001110000100011011: color_data = 12'b111011101110;
20'b01001110000100011100: color_data = 12'b111011101110;
20'b01001110000100011101: color_data = 12'b111011101110;
20'b01001110000100011110: color_data = 12'b111011101110;
20'b01001110000100011111: color_data = 12'b111011101110;
20'b01001110000100100000: color_data = 12'b111011101110;
20'b01001110000100100001: color_data = 12'b111011101110;
20'b01001110000100100010: color_data = 12'b111011101110;
20'b01001110000100100100: color_data = 12'b111011101110;
20'b01001110000100100101: color_data = 12'b111011101110;
20'b01001110000100100110: color_data = 12'b111011101110;
20'b01001110000100100111: color_data = 12'b111011101110;
20'b01001110000100101000: color_data = 12'b111011101110;
20'b01001110000100101001: color_data = 12'b111011101110;
20'b01001110000100101010: color_data = 12'b111011101110;
20'b01001110000100101011: color_data = 12'b111011101110;
20'b01001110000100101100: color_data = 12'b111011101110;
20'b01001110000100101101: color_data = 12'b111011101110;
20'b01001110000100101111: color_data = 12'b111011101110;
20'b01001110000100110000: color_data = 12'b111011101110;
20'b01001110000100110001: color_data = 12'b111011101110;
20'b01001110000100110010: color_data = 12'b111011101110;
20'b01001110000100110011: color_data = 12'b111011101110;
20'b01001110000100110100: color_data = 12'b111011101110;
20'b01001110000100110101: color_data = 12'b111011101110;
20'b01001110000100110110: color_data = 12'b111011101110;
20'b01001110000100110111: color_data = 12'b111011101110;
20'b01001110000100111000: color_data = 12'b111011101110;
20'b01001110000101000100: color_data = 12'b111011101110;
20'b01001110000101000101: color_data = 12'b111011101110;
20'b01001110000101000110: color_data = 12'b111011101110;
20'b01001110000101000111: color_data = 12'b111011101110;
20'b01001110000101001000: color_data = 12'b111011101110;
20'b01001110000101001001: color_data = 12'b111011101110;
20'b01001110000101001010: color_data = 12'b111011101110;
20'b01001110000101001011: color_data = 12'b111011101110;
20'b01001110000101001100: color_data = 12'b111011101110;
20'b01001110000101001101: color_data = 12'b111011101110;
20'b01001110000101001111: color_data = 12'b111011101110;
20'b01001110000101010000: color_data = 12'b111011101110;
20'b01001110000101010001: color_data = 12'b111011101110;
20'b01001110000101010010: color_data = 12'b111011101110;
20'b01001110000101010011: color_data = 12'b111011101110;
20'b01001110000101010100: color_data = 12'b111011101110;
20'b01001110000101010101: color_data = 12'b111011101110;
20'b01001110000101010110: color_data = 12'b111011101110;
20'b01001110000101010111: color_data = 12'b111011101110;
20'b01001110000101011000: color_data = 12'b111011101110;
20'b01001110000110011100: color_data = 12'b111011101110;
20'b01001110000110011101: color_data = 12'b111011101110;
20'b01001110000110011110: color_data = 12'b111011101110;
20'b01001110000110011111: color_data = 12'b111011101110;
20'b01001110000110100000: color_data = 12'b111011101110;
20'b01001110000110100001: color_data = 12'b111011101110;
20'b01001110000110100010: color_data = 12'b111011101110;
20'b01001110000110100011: color_data = 12'b111011101110;
20'b01001110000110100100: color_data = 12'b111011101110;
20'b01001110000110100101: color_data = 12'b111011101110;
20'b01001110000110100111: color_data = 12'b111011101110;
20'b01001110000110101000: color_data = 12'b111011101110;
20'b01001110000110101001: color_data = 12'b111011101110;
20'b01001110000110101010: color_data = 12'b111011101110;
20'b01001110000110101011: color_data = 12'b111011101110;
20'b01001110000110101100: color_data = 12'b111011101110;
20'b01001110000110101101: color_data = 12'b111011101110;
20'b01001110000110101110: color_data = 12'b111011101110;
20'b01001110000110101111: color_data = 12'b111011101110;
20'b01001110000110110000: color_data = 12'b111011101110;
20'b01001110000110111101: color_data = 12'b111011101110;
20'b01001110000110111110: color_data = 12'b111011101110;
20'b01001110000110111111: color_data = 12'b111011101110;
20'b01001110000111000000: color_data = 12'b111011101110;
20'b01001110000111000001: color_data = 12'b111011101110;
20'b01001110000111000010: color_data = 12'b111011101110;
20'b01001110000111000011: color_data = 12'b111011101110;
20'b01001110000111000100: color_data = 12'b111011101110;
20'b01001110000111000101: color_data = 12'b111011101110;
20'b01001110000111000110: color_data = 12'b111011101110;
20'b01001110000111001000: color_data = 12'b111011101110;
20'b01001110000111001001: color_data = 12'b111011101110;
20'b01001110000111001010: color_data = 12'b111011101110;
20'b01001110000111001011: color_data = 12'b111011101110;
20'b01001110000111001100: color_data = 12'b111011101110;
20'b01001110000111001101: color_data = 12'b111011101110;
20'b01001110000111001110: color_data = 12'b111011101110;
20'b01001110000111001111: color_data = 12'b111011101110;
20'b01001110000111010000: color_data = 12'b111011101110;
20'b01001110000111010001: color_data = 12'b111011101110;
20'b01001110010010010110: color_data = 12'b111011101110;
20'b01001110010010010111: color_data = 12'b111011101110;
20'b01001110010010011000: color_data = 12'b111011101110;
20'b01001110010010011001: color_data = 12'b111011101110;
20'b01001110010010011010: color_data = 12'b111011101110;
20'b01001110010010011011: color_data = 12'b111011101110;
20'b01001110010010011100: color_data = 12'b111011101110;
20'b01001110010010011101: color_data = 12'b111011101110;
20'b01001110010010011110: color_data = 12'b111011101110;
20'b01001110010010011111: color_data = 12'b111011101110;
20'b01001110010010100001: color_data = 12'b111011101110;
20'b01001110010010100010: color_data = 12'b111011101110;
20'b01001110010010100011: color_data = 12'b111011101110;
20'b01001110010010100100: color_data = 12'b111011101110;
20'b01001110010010100101: color_data = 12'b111011101110;
20'b01001110010010100110: color_data = 12'b111011101110;
20'b01001110010010100111: color_data = 12'b111011101110;
20'b01001110010010101000: color_data = 12'b111011101110;
20'b01001110010010101001: color_data = 12'b111011101110;
20'b01001110010010101010: color_data = 12'b111011101110;
20'b01001110010011001101: color_data = 12'b111011101110;
20'b01001110010011001110: color_data = 12'b111011101110;
20'b01001110010011001111: color_data = 12'b111011101110;
20'b01001110010011010000: color_data = 12'b111011101110;
20'b01001110010011010001: color_data = 12'b111011101110;
20'b01001110010011010010: color_data = 12'b111011101110;
20'b01001110010011010011: color_data = 12'b111011101110;
20'b01001110010011010100: color_data = 12'b111011101110;
20'b01001110010011010101: color_data = 12'b111011101110;
20'b01001110010011010110: color_data = 12'b111011101110;
20'b01001110010011011000: color_data = 12'b111011101110;
20'b01001110010011011001: color_data = 12'b111011101110;
20'b01001110010011011010: color_data = 12'b111011101110;
20'b01001110010011011011: color_data = 12'b111011101110;
20'b01001110010011011100: color_data = 12'b111011101110;
20'b01001110010011011101: color_data = 12'b111011101110;
20'b01001110010011011110: color_data = 12'b111011101110;
20'b01001110010011011111: color_data = 12'b111011101110;
20'b01001110010011100000: color_data = 12'b111011101110;
20'b01001110010011100001: color_data = 12'b111011101110;
20'b01001110010011101101: color_data = 12'b111011101110;
20'b01001110010011101110: color_data = 12'b111011101110;
20'b01001110010011101111: color_data = 12'b111011101110;
20'b01001110010011110000: color_data = 12'b111011101110;
20'b01001110010011110001: color_data = 12'b111011101110;
20'b01001110010011110010: color_data = 12'b111011101110;
20'b01001110010011110011: color_data = 12'b111011101110;
20'b01001110010011110100: color_data = 12'b111011101110;
20'b01001110010011110101: color_data = 12'b111011101110;
20'b01001110010011110110: color_data = 12'b111011101110;
20'b01001110010011111000: color_data = 12'b111011101110;
20'b01001110010011111001: color_data = 12'b111011101110;
20'b01001110010011111010: color_data = 12'b111011101110;
20'b01001110010011111011: color_data = 12'b111011101110;
20'b01001110010011111100: color_data = 12'b111011101110;
20'b01001110010011111101: color_data = 12'b111011101110;
20'b01001110010011111110: color_data = 12'b111011101110;
20'b01001110010011111111: color_data = 12'b111011101110;
20'b01001110010100000000: color_data = 12'b111011101110;
20'b01001110010100000001: color_data = 12'b111011101110;
20'b01001110010100000011: color_data = 12'b111011101110;
20'b01001110010100000100: color_data = 12'b111011101110;
20'b01001110010100000101: color_data = 12'b111011101110;
20'b01001110010100000110: color_data = 12'b111011101110;
20'b01001110010100000111: color_data = 12'b111011101110;
20'b01001110010100001000: color_data = 12'b111011101110;
20'b01001110010100001001: color_data = 12'b111011101110;
20'b01001110010100001010: color_data = 12'b111011101110;
20'b01001110010100001011: color_data = 12'b111011101110;
20'b01001110010100001100: color_data = 12'b111011101110;
20'b01001110010100011001: color_data = 12'b111011101110;
20'b01001110010100011010: color_data = 12'b111011101110;
20'b01001110010100011011: color_data = 12'b111011101110;
20'b01001110010100011100: color_data = 12'b111011101110;
20'b01001110010100011101: color_data = 12'b111011101110;
20'b01001110010100011110: color_data = 12'b111011101110;
20'b01001110010100011111: color_data = 12'b111011101110;
20'b01001110010100100000: color_data = 12'b111011101110;
20'b01001110010100100001: color_data = 12'b111011101110;
20'b01001110010100100010: color_data = 12'b111011101110;
20'b01001110010100100100: color_data = 12'b111011101110;
20'b01001110010100100101: color_data = 12'b111011101110;
20'b01001110010100100110: color_data = 12'b111011101110;
20'b01001110010100100111: color_data = 12'b111011101110;
20'b01001110010100101000: color_data = 12'b111011101110;
20'b01001110010100101001: color_data = 12'b111011101110;
20'b01001110010100101010: color_data = 12'b111011101110;
20'b01001110010100101011: color_data = 12'b111011101110;
20'b01001110010100101100: color_data = 12'b111011101110;
20'b01001110010100101101: color_data = 12'b111011101110;
20'b01001110010100101111: color_data = 12'b111011101110;
20'b01001110010100110000: color_data = 12'b111011101110;
20'b01001110010100110001: color_data = 12'b111011101110;
20'b01001110010100110010: color_data = 12'b111011101110;
20'b01001110010100110011: color_data = 12'b111011101110;
20'b01001110010100110100: color_data = 12'b111011101110;
20'b01001110010100110101: color_data = 12'b111011101110;
20'b01001110010100110110: color_data = 12'b111011101110;
20'b01001110010100110111: color_data = 12'b111011101110;
20'b01001110010100111000: color_data = 12'b111011101110;
20'b01001110010101000100: color_data = 12'b111011101110;
20'b01001110010101000101: color_data = 12'b111011101110;
20'b01001110010101000110: color_data = 12'b111011101110;
20'b01001110010101000111: color_data = 12'b111011101110;
20'b01001110010101001000: color_data = 12'b111011101110;
20'b01001110010101001001: color_data = 12'b111011101110;
20'b01001110010101001010: color_data = 12'b111011101110;
20'b01001110010101001011: color_data = 12'b111011101110;
20'b01001110010101001100: color_data = 12'b111011101110;
20'b01001110010101001101: color_data = 12'b111011101110;
20'b01001110010101001111: color_data = 12'b111011101110;
20'b01001110010101010000: color_data = 12'b111011101110;
20'b01001110010101010001: color_data = 12'b111011101110;
20'b01001110010101010010: color_data = 12'b111011101110;
20'b01001110010101010011: color_data = 12'b111011101110;
20'b01001110010101010100: color_data = 12'b111011101110;
20'b01001110010101010101: color_data = 12'b111011101110;
20'b01001110010101010110: color_data = 12'b111011101110;
20'b01001110010101010111: color_data = 12'b111011101110;
20'b01001110010101011000: color_data = 12'b111011101110;
20'b01001110010110011100: color_data = 12'b111011101110;
20'b01001110010110011101: color_data = 12'b111011101110;
20'b01001110010110011110: color_data = 12'b111011101110;
20'b01001110010110011111: color_data = 12'b111011101110;
20'b01001110010110100000: color_data = 12'b111011101110;
20'b01001110010110100001: color_data = 12'b111011101110;
20'b01001110010110100010: color_data = 12'b111011101110;
20'b01001110010110100011: color_data = 12'b111011101110;
20'b01001110010110100100: color_data = 12'b111011101110;
20'b01001110010110100101: color_data = 12'b111011101110;
20'b01001110010110100111: color_data = 12'b111011101110;
20'b01001110010110101000: color_data = 12'b111011101110;
20'b01001110010110101001: color_data = 12'b111011101110;
20'b01001110010110101010: color_data = 12'b111011101110;
20'b01001110010110101011: color_data = 12'b111011101110;
20'b01001110010110101100: color_data = 12'b111011101110;
20'b01001110010110101101: color_data = 12'b111011101110;
20'b01001110010110101110: color_data = 12'b111011101110;
20'b01001110010110101111: color_data = 12'b111011101110;
20'b01001110010110110000: color_data = 12'b111011101110;
20'b01001110010110111101: color_data = 12'b111011101110;
20'b01001110010110111110: color_data = 12'b111011101110;
20'b01001110010110111111: color_data = 12'b111011101110;
20'b01001110010111000000: color_data = 12'b111011101110;
20'b01001110010111000001: color_data = 12'b111011101110;
20'b01001110010111000010: color_data = 12'b111011101110;
20'b01001110010111000011: color_data = 12'b111011101110;
20'b01001110010111000100: color_data = 12'b111011101110;
20'b01001110010111000101: color_data = 12'b111011101110;
20'b01001110010111000110: color_data = 12'b111011101110;
20'b01001110010111001000: color_data = 12'b111011101110;
20'b01001110010111001001: color_data = 12'b111011101110;
20'b01001110010111001010: color_data = 12'b111011101110;
20'b01001110010111001011: color_data = 12'b111011101110;
20'b01001110010111001100: color_data = 12'b111011101110;
20'b01001110010111001101: color_data = 12'b111011101110;
20'b01001110010111001110: color_data = 12'b111011101110;
20'b01001110010111001111: color_data = 12'b111011101110;
20'b01001110010111010000: color_data = 12'b111011101110;
20'b01001110010111010001: color_data = 12'b111011101110;
20'b01001110100010010110: color_data = 12'b111011101110;
20'b01001110100010010111: color_data = 12'b111011101110;
20'b01001110100010011000: color_data = 12'b111011101110;
20'b01001110100010011001: color_data = 12'b111011101110;
20'b01001110100010011010: color_data = 12'b111011101110;
20'b01001110100010011011: color_data = 12'b111011101110;
20'b01001110100010011100: color_data = 12'b111011101110;
20'b01001110100010011101: color_data = 12'b111011101110;
20'b01001110100010011110: color_data = 12'b111011101110;
20'b01001110100010011111: color_data = 12'b111011101110;
20'b01001110100010100001: color_data = 12'b111011101110;
20'b01001110100010100010: color_data = 12'b111011101110;
20'b01001110100010100011: color_data = 12'b111011101110;
20'b01001110100010100100: color_data = 12'b111011101110;
20'b01001110100010100101: color_data = 12'b111011101110;
20'b01001110100010100110: color_data = 12'b111011101110;
20'b01001110100010100111: color_data = 12'b111011101110;
20'b01001110100010101000: color_data = 12'b111011101110;
20'b01001110100010101001: color_data = 12'b111011101110;
20'b01001110100010101010: color_data = 12'b111011101110;
20'b01001110100011001101: color_data = 12'b111011101110;
20'b01001110100011001110: color_data = 12'b111011101110;
20'b01001110100011001111: color_data = 12'b111011101110;
20'b01001110100011010000: color_data = 12'b111011101110;
20'b01001110100011010001: color_data = 12'b111011101110;
20'b01001110100011010010: color_data = 12'b111011101110;
20'b01001110100011010011: color_data = 12'b111011101110;
20'b01001110100011010100: color_data = 12'b111011101110;
20'b01001110100011010101: color_data = 12'b111011101110;
20'b01001110100011010110: color_data = 12'b111011101110;
20'b01001110100011011000: color_data = 12'b111011101110;
20'b01001110100011011001: color_data = 12'b111011101110;
20'b01001110100011011010: color_data = 12'b111011101110;
20'b01001110100011011011: color_data = 12'b111011101110;
20'b01001110100011011100: color_data = 12'b111011101110;
20'b01001110100011011101: color_data = 12'b111011101110;
20'b01001110100011011110: color_data = 12'b111011101110;
20'b01001110100011011111: color_data = 12'b111011101110;
20'b01001110100011100000: color_data = 12'b111011101110;
20'b01001110100011100001: color_data = 12'b111011101110;
20'b01001110100011101101: color_data = 12'b111011101110;
20'b01001110100011101110: color_data = 12'b111011101110;
20'b01001110100011101111: color_data = 12'b111011101110;
20'b01001110100011110000: color_data = 12'b111011101110;
20'b01001110100011110001: color_data = 12'b111011101110;
20'b01001110100011110010: color_data = 12'b111011101110;
20'b01001110100011110011: color_data = 12'b111011101110;
20'b01001110100011110100: color_data = 12'b111011101110;
20'b01001110100011110101: color_data = 12'b111011101110;
20'b01001110100011110110: color_data = 12'b111011101110;
20'b01001110100011111000: color_data = 12'b111011101110;
20'b01001110100011111001: color_data = 12'b111011101110;
20'b01001110100011111010: color_data = 12'b111011101110;
20'b01001110100011111011: color_data = 12'b111011101110;
20'b01001110100011111100: color_data = 12'b111011101110;
20'b01001110100011111101: color_data = 12'b111011101110;
20'b01001110100011111110: color_data = 12'b111011101110;
20'b01001110100011111111: color_data = 12'b111011101110;
20'b01001110100100000000: color_data = 12'b111011101110;
20'b01001110100100000001: color_data = 12'b111011101110;
20'b01001110100100000011: color_data = 12'b111011101110;
20'b01001110100100000100: color_data = 12'b111011101110;
20'b01001110100100000101: color_data = 12'b111011101110;
20'b01001110100100000110: color_data = 12'b111011101110;
20'b01001110100100000111: color_data = 12'b111011101110;
20'b01001110100100001000: color_data = 12'b111011101110;
20'b01001110100100001001: color_data = 12'b111011101110;
20'b01001110100100001010: color_data = 12'b111011101110;
20'b01001110100100001011: color_data = 12'b111011101110;
20'b01001110100100001100: color_data = 12'b111011101110;
20'b01001110100100011001: color_data = 12'b111011101110;
20'b01001110100100011010: color_data = 12'b111011101110;
20'b01001110100100011011: color_data = 12'b111011101110;
20'b01001110100100011100: color_data = 12'b111011101110;
20'b01001110100100011101: color_data = 12'b111011101110;
20'b01001110100100011110: color_data = 12'b111011101110;
20'b01001110100100011111: color_data = 12'b111011101110;
20'b01001110100100100000: color_data = 12'b111011101110;
20'b01001110100100100001: color_data = 12'b111011101110;
20'b01001110100100100010: color_data = 12'b111011101110;
20'b01001110100100100100: color_data = 12'b111011101110;
20'b01001110100100100101: color_data = 12'b111011101110;
20'b01001110100100100110: color_data = 12'b111011101110;
20'b01001110100100100111: color_data = 12'b111011101110;
20'b01001110100100101000: color_data = 12'b111011101110;
20'b01001110100100101001: color_data = 12'b111011101110;
20'b01001110100100101010: color_data = 12'b111011101110;
20'b01001110100100101011: color_data = 12'b111011101110;
20'b01001110100100101100: color_data = 12'b111011101110;
20'b01001110100100101101: color_data = 12'b111011101110;
20'b01001110100100101111: color_data = 12'b111011101110;
20'b01001110100100110000: color_data = 12'b111011101110;
20'b01001110100100110001: color_data = 12'b111011101110;
20'b01001110100100110010: color_data = 12'b111011101110;
20'b01001110100100110011: color_data = 12'b111011101110;
20'b01001110100100110100: color_data = 12'b111011101110;
20'b01001110100100110101: color_data = 12'b111011101110;
20'b01001110100100110110: color_data = 12'b111011101110;
20'b01001110100100110111: color_data = 12'b111011101110;
20'b01001110100100111000: color_data = 12'b111011101110;
20'b01001110100101000100: color_data = 12'b111011101110;
20'b01001110100101000101: color_data = 12'b111011101110;
20'b01001110100101000110: color_data = 12'b111011101110;
20'b01001110100101000111: color_data = 12'b111011101110;
20'b01001110100101001000: color_data = 12'b111011101110;
20'b01001110100101001001: color_data = 12'b111011101110;
20'b01001110100101001010: color_data = 12'b111011101110;
20'b01001110100101001011: color_data = 12'b111011101110;
20'b01001110100101001100: color_data = 12'b111011101110;
20'b01001110100101001101: color_data = 12'b111011101110;
20'b01001110100101001111: color_data = 12'b111011101110;
20'b01001110100101010000: color_data = 12'b111011101110;
20'b01001110100101010001: color_data = 12'b111011101110;
20'b01001110100101010010: color_data = 12'b111011101110;
20'b01001110100101010011: color_data = 12'b111011101110;
20'b01001110100101010100: color_data = 12'b111011101110;
20'b01001110100101010101: color_data = 12'b111011101110;
20'b01001110100101010110: color_data = 12'b111011101110;
20'b01001110100101010111: color_data = 12'b111011101110;
20'b01001110100101011000: color_data = 12'b111011101110;
20'b01001110100110011100: color_data = 12'b111011101110;
20'b01001110100110011101: color_data = 12'b111011101110;
20'b01001110100110011110: color_data = 12'b111011101110;
20'b01001110100110011111: color_data = 12'b111011101110;
20'b01001110100110100000: color_data = 12'b111011101110;
20'b01001110100110100001: color_data = 12'b111011101110;
20'b01001110100110100010: color_data = 12'b111011101110;
20'b01001110100110100011: color_data = 12'b111011101110;
20'b01001110100110100100: color_data = 12'b111011101110;
20'b01001110100110100101: color_data = 12'b111011101110;
20'b01001110100110100111: color_data = 12'b111011101110;
20'b01001110100110101000: color_data = 12'b111011101110;
20'b01001110100110101001: color_data = 12'b111011101110;
20'b01001110100110101010: color_data = 12'b111011101110;
20'b01001110100110101011: color_data = 12'b111011101110;
20'b01001110100110101100: color_data = 12'b111011101110;
20'b01001110100110101101: color_data = 12'b111011101110;
20'b01001110100110101110: color_data = 12'b111011101110;
20'b01001110100110101111: color_data = 12'b111011101110;
20'b01001110100110110000: color_data = 12'b111011101110;
20'b01001110100110111101: color_data = 12'b111011101110;
20'b01001110100110111110: color_data = 12'b111011101110;
20'b01001110100110111111: color_data = 12'b111011101110;
20'b01001110100111000000: color_data = 12'b111011101110;
20'b01001110100111000001: color_data = 12'b111011101110;
20'b01001110100111000010: color_data = 12'b111011101110;
20'b01001110100111000011: color_data = 12'b111011101110;
20'b01001110100111000100: color_data = 12'b111011101110;
20'b01001110100111000101: color_data = 12'b111011101110;
20'b01001110100111000110: color_data = 12'b111011101110;
20'b01001110100111001000: color_data = 12'b111011101110;
20'b01001110100111001001: color_data = 12'b111011101110;
20'b01001110100111001010: color_data = 12'b111011101110;
20'b01001110100111001011: color_data = 12'b111011101110;
20'b01001110100111001100: color_data = 12'b111011101110;
20'b01001110100111001101: color_data = 12'b111011101110;
20'b01001110100111001110: color_data = 12'b111011101110;
20'b01001110100111001111: color_data = 12'b111011101110;
20'b01001110100111010000: color_data = 12'b111011101110;
20'b01001110100111010001: color_data = 12'b111011101110;
20'b01001110110010010110: color_data = 12'b111011101110;
20'b01001110110010010111: color_data = 12'b111011101110;
20'b01001110110010011000: color_data = 12'b111011101110;
20'b01001110110010011001: color_data = 12'b111011101110;
20'b01001110110010011010: color_data = 12'b111011101110;
20'b01001110110010011011: color_data = 12'b111011101110;
20'b01001110110010011100: color_data = 12'b111011101110;
20'b01001110110010011101: color_data = 12'b111011101110;
20'b01001110110010011110: color_data = 12'b111011101110;
20'b01001110110010011111: color_data = 12'b111011101110;
20'b01001110110010100001: color_data = 12'b111011101110;
20'b01001110110010100010: color_data = 12'b111011101110;
20'b01001110110010100011: color_data = 12'b111011101110;
20'b01001110110010100100: color_data = 12'b111011101110;
20'b01001110110010100101: color_data = 12'b111011101110;
20'b01001110110010100110: color_data = 12'b111011101110;
20'b01001110110010100111: color_data = 12'b111011101110;
20'b01001110110010101000: color_data = 12'b111011101110;
20'b01001110110010101001: color_data = 12'b111011101110;
20'b01001110110010101010: color_data = 12'b111011101110;
20'b01001110110011001101: color_data = 12'b111011101110;
20'b01001110110011001110: color_data = 12'b111011101110;
20'b01001110110011001111: color_data = 12'b111011101110;
20'b01001110110011010000: color_data = 12'b111011101110;
20'b01001110110011010001: color_data = 12'b111011101110;
20'b01001110110011010010: color_data = 12'b111011101110;
20'b01001110110011010011: color_data = 12'b111011101110;
20'b01001110110011010100: color_data = 12'b111011101110;
20'b01001110110011010101: color_data = 12'b111011101110;
20'b01001110110011010110: color_data = 12'b111011101110;
20'b01001110110011011000: color_data = 12'b111011101110;
20'b01001110110011011001: color_data = 12'b111011101110;
20'b01001110110011011010: color_data = 12'b111011101110;
20'b01001110110011011011: color_data = 12'b111011101110;
20'b01001110110011011100: color_data = 12'b111011101110;
20'b01001110110011011101: color_data = 12'b111011101110;
20'b01001110110011011110: color_data = 12'b111011101110;
20'b01001110110011011111: color_data = 12'b111011101110;
20'b01001110110011100000: color_data = 12'b111011101110;
20'b01001110110011100001: color_data = 12'b111011101110;
20'b01001110110011101101: color_data = 12'b111011101110;
20'b01001110110011101110: color_data = 12'b111011101110;
20'b01001110110011101111: color_data = 12'b111011101110;
20'b01001110110011110000: color_data = 12'b111011101110;
20'b01001110110011110001: color_data = 12'b111011101110;
20'b01001110110011110010: color_data = 12'b111011101110;
20'b01001110110011110011: color_data = 12'b111011101110;
20'b01001110110011110100: color_data = 12'b111011101110;
20'b01001110110011110101: color_data = 12'b111011101110;
20'b01001110110011110110: color_data = 12'b111011101110;
20'b01001110110011111000: color_data = 12'b111011101110;
20'b01001110110011111001: color_data = 12'b111011101110;
20'b01001110110011111010: color_data = 12'b111011101110;
20'b01001110110011111011: color_data = 12'b111011101110;
20'b01001110110011111100: color_data = 12'b111011101110;
20'b01001110110011111101: color_data = 12'b111011101110;
20'b01001110110011111110: color_data = 12'b111011101110;
20'b01001110110011111111: color_data = 12'b111011101110;
20'b01001110110100000000: color_data = 12'b111011101110;
20'b01001110110100000001: color_data = 12'b111011101110;
20'b01001110110100000011: color_data = 12'b111011101110;
20'b01001110110100000100: color_data = 12'b111011101110;
20'b01001110110100000101: color_data = 12'b111011101110;
20'b01001110110100000110: color_data = 12'b111011101110;
20'b01001110110100000111: color_data = 12'b111011101110;
20'b01001110110100001000: color_data = 12'b111011101110;
20'b01001110110100001001: color_data = 12'b111011101110;
20'b01001110110100001010: color_data = 12'b111011101110;
20'b01001110110100001011: color_data = 12'b111011101110;
20'b01001110110100001100: color_data = 12'b111011101110;
20'b01001110110100011001: color_data = 12'b111011101110;
20'b01001110110100011010: color_data = 12'b111011101110;
20'b01001110110100011011: color_data = 12'b111011101110;
20'b01001110110100011100: color_data = 12'b111011101110;
20'b01001110110100011101: color_data = 12'b111011101110;
20'b01001110110100011110: color_data = 12'b111011101110;
20'b01001110110100011111: color_data = 12'b111011101110;
20'b01001110110100100000: color_data = 12'b111011101110;
20'b01001110110100100001: color_data = 12'b111011101110;
20'b01001110110100100010: color_data = 12'b111011101110;
20'b01001110110100100100: color_data = 12'b111011101110;
20'b01001110110100100101: color_data = 12'b111011101110;
20'b01001110110100100110: color_data = 12'b111011101110;
20'b01001110110100100111: color_data = 12'b111011101110;
20'b01001110110100101000: color_data = 12'b111011101110;
20'b01001110110100101001: color_data = 12'b111011101110;
20'b01001110110100101010: color_data = 12'b111011101110;
20'b01001110110100101011: color_data = 12'b111011101110;
20'b01001110110100101100: color_data = 12'b111011101110;
20'b01001110110100101101: color_data = 12'b111011101110;
20'b01001110110100101111: color_data = 12'b111011101110;
20'b01001110110100110000: color_data = 12'b111011101110;
20'b01001110110100110001: color_data = 12'b111011101110;
20'b01001110110100110010: color_data = 12'b111011101110;
20'b01001110110100110011: color_data = 12'b111011101110;
20'b01001110110100110100: color_data = 12'b111011101110;
20'b01001110110100110101: color_data = 12'b111011101110;
20'b01001110110100110110: color_data = 12'b111011101110;
20'b01001110110100110111: color_data = 12'b111011101110;
20'b01001110110100111000: color_data = 12'b111011101110;
20'b01001110110101000100: color_data = 12'b111011101110;
20'b01001110110101000101: color_data = 12'b111011101110;
20'b01001110110101000110: color_data = 12'b111011101110;
20'b01001110110101000111: color_data = 12'b111011101110;
20'b01001110110101001000: color_data = 12'b111011101110;
20'b01001110110101001001: color_data = 12'b111011101110;
20'b01001110110101001010: color_data = 12'b111011101110;
20'b01001110110101001011: color_data = 12'b111011101110;
20'b01001110110101001100: color_data = 12'b111011101110;
20'b01001110110101001101: color_data = 12'b111011101110;
20'b01001110110101001111: color_data = 12'b111011101110;
20'b01001110110101010000: color_data = 12'b111011101110;
20'b01001110110101010001: color_data = 12'b111011101110;
20'b01001110110101010010: color_data = 12'b111011101110;
20'b01001110110101010011: color_data = 12'b111011101110;
20'b01001110110101010100: color_data = 12'b111011101110;
20'b01001110110101010101: color_data = 12'b111011101110;
20'b01001110110101010110: color_data = 12'b111011101110;
20'b01001110110101010111: color_data = 12'b111011101110;
20'b01001110110101011000: color_data = 12'b111011101110;
20'b01001110110110011100: color_data = 12'b111011101110;
20'b01001110110110011101: color_data = 12'b111011101110;
20'b01001110110110011110: color_data = 12'b111011101110;
20'b01001110110110011111: color_data = 12'b111011101110;
20'b01001110110110100000: color_data = 12'b111011101110;
20'b01001110110110100001: color_data = 12'b111011101110;
20'b01001110110110100010: color_data = 12'b111011101110;
20'b01001110110110100011: color_data = 12'b111011101110;
20'b01001110110110100100: color_data = 12'b111011101110;
20'b01001110110110100101: color_data = 12'b111011101110;
20'b01001110110110100111: color_data = 12'b111011101110;
20'b01001110110110101000: color_data = 12'b111011101110;
20'b01001110110110101001: color_data = 12'b111011101110;
20'b01001110110110101010: color_data = 12'b111011101110;
20'b01001110110110101011: color_data = 12'b111011101110;
20'b01001110110110101100: color_data = 12'b111011101110;
20'b01001110110110101101: color_data = 12'b111011101110;
20'b01001110110110101110: color_data = 12'b111011101110;
20'b01001110110110101111: color_data = 12'b111011101110;
20'b01001110110110110000: color_data = 12'b111011101110;
20'b01001110110110111101: color_data = 12'b111011101110;
20'b01001110110110111110: color_data = 12'b111011101110;
20'b01001110110110111111: color_data = 12'b111011101110;
20'b01001110110111000000: color_data = 12'b111011101110;
20'b01001110110111000001: color_data = 12'b111011101110;
20'b01001110110111000010: color_data = 12'b111011101110;
20'b01001110110111000011: color_data = 12'b111011101110;
20'b01001110110111000100: color_data = 12'b111011101110;
20'b01001110110111000101: color_data = 12'b111011101110;
20'b01001110110111000110: color_data = 12'b111011101110;
20'b01001110110111001000: color_data = 12'b111011101110;
20'b01001110110111001001: color_data = 12'b111011101110;
20'b01001110110111001010: color_data = 12'b111011101110;
20'b01001110110111001011: color_data = 12'b111011101110;
20'b01001110110111001100: color_data = 12'b111011101110;
20'b01001110110111001101: color_data = 12'b111011101110;
20'b01001110110111001110: color_data = 12'b111011101110;
20'b01001110110111001111: color_data = 12'b111011101110;
20'b01001110110111010000: color_data = 12'b111011101110;
20'b01001110110111010001: color_data = 12'b111011101110;
20'b01001111000010010110: color_data = 12'b111011101110;
20'b01001111000010010111: color_data = 12'b111011101110;
20'b01001111000010011000: color_data = 12'b111011101110;
20'b01001111000010011001: color_data = 12'b111011101110;
20'b01001111000010011010: color_data = 12'b111011101110;
20'b01001111000010011011: color_data = 12'b111011101110;
20'b01001111000010011100: color_data = 12'b111011101110;
20'b01001111000010011101: color_data = 12'b111011101110;
20'b01001111000010011110: color_data = 12'b111011101110;
20'b01001111000010011111: color_data = 12'b111011101110;
20'b01001111000010100001: color_data = 12'b111011101110;
20'b01001111000010100010: color_data = 12'b111011101110;
20'b01001111000010100011: color_data = 12'b111011101110;
20'b01001111000010100100: color_data = 12'b111011101110;
20'b01001111000010100101: color_data = 12'b111011101110;
20'b01001111000010100110: color_data = 12'b111011101110;
20'b01001111000010100111: color_data = 12'b111011101110;
20'b01001111000010101000: color_data = 12'b111011101110;
20'b01001111000010101001: color_data = 12'b111011101110;
20'b01001111000010101010: color_data = 12'b111011101110;
20'b01001111000011001101: color_data = 12'b111011101110;
20'b01001111000011001110: color_data = 12'b111011101110;
20'b01001111000011001111: color_data = 12'b111011101110;
20'b01001111000011010000: color_data = 12'b111011101110;
20'b01001111000011010001: color_data = 12'b111011101110;
20'b01001111000011010010: color_data = 12'b111011101110;
20'b01001111000011010011: color_data = 12'b111011101110;
20'b01001111000011010100: color_data = 12'b111011101110;
20'b01001111000011010101: color_data = 12'b111011101110;
20'b01001111000011010110: color_data = 12'b111011101110;
20'b01001111000011011000: color_data = 12'b111011101110;
20'b01001111000011011001: color_data = 12'b111011101110;
20'b01001111000011011010: color_data = 12'b111011101110;
20'b01001111000011011011: color_data = 12'b111011101110;
20'b01001111000011011100: color_data = 12'b111011101110;
20'b01001111000011011101: color_data = 12'b111011101110;
20'b01001111000011011110: color_data = 12'b111011101110;
20'b01001111000011011111: color_data = 12'b111011101110;
20'b01001111000011100000: color_data = 12'b111011101110;
20'b01001111000011100001: color_data = 12'b111011101110;
20'b01001111000011101101: color_data = 12'b111011101110;
20'b01001111000011101110: color_data = 12'b111011101110;
20'b01001111000011101111: color_data = 12'b111011101110;
20'b01001111000011110000: color_data = 12'b111011101110;
20'b01001111000011110001: color_data = 12'b111011101110;
20'b01001111000011110010: color_data = 12'b111011101110;
20'b01001111000011110011: color_data = 12'b111011101110;
20'b01001111000011110100: color_data = 12'b111011101110;
20'b01001111000011110101: color_data = 12'b111011101110;
20'b01001111000011110110: color_data = 12'b111011101110;
20'b01001111000011111000: color_data = 12'b111011101110;
20'b01001111000011111001: color_data = 12'b111011101110;
20'b01001111000011111010: color_data = 12'b111011101110;
20'b01001111000011111011: color_data = 12'b111011101110;
20'b01001111000011111100: color_data = 12'b111011101110;
20'b01001111000011111101: color_data = 12'b111011101110;
20'b01001111000011111110: color_data = 12'b111011101110;
20'b01001111000011111111: color_data = 12'b111011101110;
20'b01001111000100000000: color_data = 12'b111011101110;
20'b01001111000100000001: color_data = 12'b111011101110;
20'b01001111000100000011: color_data = 12'b111011101110;
20'b01001111000100000100: color_data = 12'b111011101110;
20'b01001111000100000101: color_data = 12'b111011101110;
20'b01001111000100000110: color_data = 12'b111011101110;
20'b01001111000100000111: color_data = 12'b111011101110;
20'b01001111000100001000: color_data = 12'b111011101110;
20'b01001111000100001001: color_data = 12'b111011101110;
20'b01001111000100001010: color_data = 12'b111011101110;
20'b01001111000100001011: color_data = 12'b111011101110;
20'b01001111000100001100: color_data = 12'b111011101110;
20'b01001111000100011001: color_data = 12'b111011101110;
20'b01001111000100011010: color_data = 12'b111011101110;
20'b01001111000100011011: color_data = 12'b111011101110;
20'b01001111000100011100: color_data = 12'b111011101110;
20'b01001111000100011101: color_data = 12'b111011101110;
20'b01001111000100011110: color_data = 12'b111011101110;
20'b01001111000100011111: color_data = 12'b111011101110;
20'b01001111000100100000: color_data = 12'b111011101110;
20'b01001111000100100001: color_data = 12'b111011101110;
20'b01001111000100100010: color_data = 12'b111011101110;
20'b01001111000100100100: color_data = 12'b111011101110;
20'b01001111000100100101: color_data = 12'b111011101110;
20'b01001111000100100110: color_data = 12'b111011101110;
20'b01001111000100100111: color_data = 12'b111011101110;
20'b01001111000100101000: color_data = 12'b111011101110;
20'b01001111000100101001: color_data = 12'b111011101110;
20'b01001111000100101010: color_data = 12'b111011101110;
20'b01001111000100101011: color_data = 12'b111011101110;
20'b01001111000100101100: color_data = 12'b111011101110;
20'b01001111000100101101: color_data = 12'b111011101110;
20'b01001111000100101111: color_data = 12'b111011101110;
20'b01001111000100110000: color_data = 12'b111011101110;
20'b01001111000100110001: color_data = 12'b111011101110;
20'b01001111000100110010: color_data = 12'b111011101110;
20'b01001111000100110011: color_data = 12'b111011101110;
20'b01001111000100110100: color_data = 12'b111011101110;
20'b01001111000100110101: color_data = 12'b111011101110;
20'b01001111000100110110: color_data = 12'b111011101110;
20'b01001111000100110111: color_data = 12'b111011101110;
20'b01001111000100111000: color_data = 12'b111011101110;
20'b01001111000101000100: color_data = 12'b111011101110;
20'b01001111000101000101: color_data = 12'b111011101110;
20'b01001111000101000110: color_data = 12'b111011101110;
20'b01001111000101000111: color_data = 12'b111011101110;
20'b01001111000101001000: color_data = 12'b111011101110;
20'b01001111000101001001: color_data = 12'b111011101110;
20'b01001111000101001010: color_data = 12'b111011101110;
20'b01001111000101001011: color_data = 12'b111011101110;
20'b01001111000101001100: color_data = 12'b111011101110;
20'b01001111000101001101: color_data = 12'b111011101110;
20'b01001111000101001111: color_data = 12'b111011101110;
20'b01001111000101010000: color_data = 12'b111011101110;
20'b01001111000101010001: color_data = 12'b111011101110;
20'b01001111000101010010: color_data = 12'b111011101110;
20'b01001111000101010011: color_data = 12'b111011101110;
20'b01001111000101010100: color_data = 12'b111011101110;
20'b01001111000101010101: color_data = 12'b111011101110;
20'b01001111000101010110: color_data = 12'b111011101110;
20'b01001111000101010111: color_data = 12'b111011101110;
20'b01001111000101011000: color_data = 12'b111011101110;
20'b01001111000110011100: color_data = 12'b111011101110;
20'b01001111000110011101: color_data = 12'b111011101110;
20'b01001111000110011110: color_data = 12'b111011101110;
20'b01001111000110011111: color_data = 12'b111011101110;
20'b01001111000110100000: color_data = 12'b111011101110;
20'b01001111000110100001: color_data = 12'b111011101110;
20'b01001111000110100010: color_data = 12'b111011101110;
20'b01001111000110100011: color_data = 12'b111011101110;
20'b01001111000110100100: color_data = 12'b111011101110;
20'b01001111000110100101: color_data = 12'b111011101110;
20'b01001111000110100111: color_data = 12'b111011101110;
20'b01001111000110101000: color_data = 12'b111011101110;
20'b01001111000110101001: color_data = 12'b111011101110;
20'b01001111000110101010: color_data = 12'b111011101110;
20'b01001111000110101011: color_data = 12'b111011101110;
20'b01001111000110101100: color_data = 12'b111011101110;
20'b01001111000110101101: color_data = 12'b111011101110;
20'b01001111000110101110: color_data = 12'b111011101110;
20'b01001111000110101111: color_data = 12'b111011101110;
20'b01001111000110110000: color_data = 12'b111011101110;
20'b01001111000110111101: color_data = 12'b111011101110;
20'b01001111000110111110: color_data = 12'b111011101110;
20'b01001111000110111111: color_data = 12'b111011101110;
20'b01001111000111000000: color_data = 12'b111011101110;
20'b01001111000111000001: color_data = 12'b111011101110;
20'b01001111000111000010: color_data = 12'b111011101110;
20'b01001111000111000011: color_data = 12'b111011101110;
20'b01001111000111000100: color_data = 12'b111011101110;
20'b01001111000111000101: color_data = 12'b111011101110;
20'b01001111000111000110: color_data = 12'b111011101110;
20'b01001111000111001000: color_data = 12'b111011101110;
20'b01001111000111001001: color_data = 12'b111011101110;
20'b01001111000111001010: color_data = 12'b111011101110;
20'b01001111000111001011: color_data = 12'b111011101110;
20'b01001111000111001100: color_data = 12'b111011101110;
20'b01001111000111001101: color_data = 12'b111011101110;
20'b01001111000111001110: color_data = 12'b111011101110;
20'b01001111000111001111: color_data = 12'b111011101110;
20'b01001111000111010000: color_data = 12'b111011101110;
20'b01001111000111010001: color_data = 12'b111011101110;
20'b01001111010010010110: color_data = 12'b111011101110;
20'b01001111010010010111: color_data = 12'b111011101110;
20'b01001111010010011000: color_data = 12'b111011101110;
20'b01001111010010011001: color_data = 12'b111011101110;
20'b01001111010010011010: color_data = 12'b111011101110;
20'b01001111010010011011: color_data = 12'b111011101110;
20'b01001111010010011100: color_data = 12'b111011101110;
20'b01001111010010011101: color_data = 12'b111011101110;
20'b01001111010010011110: color_data = 12'b111011101110;
20'b01001111010010011111: color_data = 12'b111011101110;
20'b01001111010010100001: color_data = 12'b111011101110;
20'b01001111010010100010: color_data = 12'b111011101110;
20'b01001111010010100011: color_data = 12'b111011101110;
20'b01001111010010100100: color_data = 12'b111011101110;
20'b01001111010010100101: color_data = 12'b111011101110;
20'b01001111010010100110: color_data = 12'b111011101110;
20'b01001111010010100111: color_data = 12'b111011101110;
20'b01001111010010101000: color_data = 12'b111011101110;
20'b01001111010010101001: color_data = 12'b111011101110;
20'b01001111010010101010: color_data = 12'b111011101110;
20'b01001111010011001101: color_data = 12'b111011101110;
20'b01001111010011001110: color_data = 12'b111011101110;
20'b01001111010011001111: color_data = 12'b111011101110;
20'b01001111010011010000: color_data = 12'b111011101110;
20'b01001111010011010001: color_data = 12'b111011101110;
20'b01001111010011010010: color_data = 12'b111011101110;
20'b01001111010011010011: color_data = 12'b111011101110;
20'b01001111010011010100: color_data = 12'b111011101110;
20'b01001111010011010101: color_data = 12'b111011101110;
20'b01001111010011010110: color_data = 12'b111011101110;
20'b01001111010011011000: color_data = 12'b111011101110;
20'b01001111010011011001: color_data = 12'b111011101110;
20'b01001111010011011010: color_data = 12'b111011101110;
20'b01001111010011011011: color_data = 12'b111011101110;
20'b01001111010011011100: color_data = 12'b111011101110;
20'b01001111010011011101: color_data = 12'b111011101110;
20'b01001111010011011110: color_data = 12'b111011101110;
20'b01001111010011011111: color_data = 12'b111011101110;
20'b01001111010011100000: color_data = 12'b111011101110;
20'b01001111010011100001: color_data = 12'b111011101110;
20'b01001111010011101101: color_data = 12'b111011101110;
20'b01001111010011101110: color_data = 12'b111011101110;
20'b01001111010011101111: color_data = 12'b111011101110;
20'b01001111010011110000: color_data = 12'b111011101110;
20'b01001111010011110001: color_data = 12'b111011101110;
20'b01001111010011110010: color_data = 12'b111011101110;
20'b01001111010011110011: color_data = 12'b111011101110;
20'b01001111010011110100: color_data = 12'b111011101110;
20'b01001111010011110101: color_data = 12'b111011101110;
20'b01001111010011110110: color_data = 12'b111011101110;
20'b01001111010011111000: color_data = 12'b111011101110;
20'b01001111010011111001: color_data = 12'b111011101110;
20'b01001111010011111010: color_data = 12'b111011101110;
20'b01001111010011111011: color_data = 12'b111011101110;
20'b01001111010011111100: color_data = 12'b111011101110;
20'b01001111010011111101: color_data = 12'b111011101110;
20'b01001111010011111110: color_data = 12'b111011101110;
20'b01001111010011111111: color_data = 12'b111011101110;
20'b01001111010100000000: color_data = 12'b111011101110;
20'b01001111010100000001: color_data = 12'b111011101110;
20'b01001111010100000011: color_data = 12'b111011101110;
20'b01001111010100000100: color_data = 12'b111011101110;
20'b01001111010100000101: color_data = 12'b111011101110;
20'b01001111010100000110: color_data = 12'b111011101110;
20'b01001111010100000111: color_data = 12'b111011101110;
20'b01001111010100001000: color_data = 12'b111011101110;
20'b01001111010100001001: color_data = 12'b111011101110;
20'b01001111010100001010: color_data = 12'b111011101110;
20'b01001111010100001011: color_data = 12'b111011101110;
20'b01001111010100001100: color_data = 12'b111011101110;
20'b01001111010100011001: color_data = 12'b111011101110;
20'b01001111010100011010: color_data = 12'b111011101110;
20'b01001111010100011011: color_data = 12'b111011101110;
20'b01001111010100011100: color_data = 12'b111011101110;
20'b01001111010100011101: color_data = 12'b111011101110;
20'b01001111010100011110: color_data = 12'b111011101110;
20'b01001111010100011111: color_data = 12'b111011101110;
20'b01001111010100100000: color_data = 12'b111011101110;
20'b01001111010100100001: color_data = 12'b111011101110;
20'b01001111010100100010: color_data = 12'b111011101110;
20'b01001111010100100100: color_data = 12'b111011101110;
20'b01001111010100100101: color_data = 12'b111011101110;
20'b01001111010100100110: color_data = 12'b111011101110;
20'b01001111010100100111: color_data = 12'b111011101110;
20'b01001111010100101000: color_data = 12'b111011101110;
20'b01001111010100101001: color_data = 12'b111011101110;
20'b01001111010100101010: color_data = 12'b111011101110;
20'b01001111010100101011: color_data = 12'b111011101110;
20'b01001111010100101100: color_data = 12'b111011101110;
20'b01001111010100101101: color_data = 12'b111011101110;
20'b01001111010100101111: color_data = 12'b111011101110;
20'b01001111010100110000: color_data = 12'b111011101110;
20'b01001111010100110001: color_data = 12'b111011101110;
20'b01001111010100110010: color_data = 12'b111011101110;
20'b01001111010100110011: color_data = 12'b111011101110;
20'b01001111010100110100: color_data = 12'b111011101110;
20'b01001111010100110101: color_data = 12'b111011101110;
20'b01001111010100110110: color_data = 12'b111011101110;
20'b01001111010100110111: color_data = 12'b111011101110;
20'b01001111010100111000: color_data = 12'b111011101110;
20'b01001111010101000100: color_data = 12'b111011101110;
20'b01001111010101000101: color_data = 12'b111011101110;
20'b01001111010101000110: color_data = 12'b111011101110;
20'b01001111010101000111: color_data = 12'b111011101110;
20'b01001111010101001000: color_data = 12'b111011101110;
20'b01001111010101001001: color_data = 12'b111011101110;
20'b01001111010101001010: color_data = 12'b111011101110;
20'b01001111010101001011: color_data = 12'b111011101110;
20'b01001111010101001100: color_data = 12'b111011101110;
20'b01001111010101001101: color_data = 12'b111011101110;
20'b01001111010101001111: color_data = 12'b111011101110;
20'b01001111010101010000: color_data = 12'b111011101110;
20'b01001111010101010001: color_data = 12'b111011101110;
20'b01001111010101010010: color_data = 12'b111011101110;
20'b01001111010101010011: color_data = 12'b111011101110;
20'b01001111010101010100: color_data = 12'b111011101110;
20'b01001111010101010101: color_data = 12'b111011101110;
20'b01001111010101010110: color_data = 12'b111011101110;
20'b01001111010101010111: color_data = 12'b111011101110;
20'b01001111010101011000: color_data = 12'b111011101110;
20'b01001111010110011100: color_data = 12'b111011101110;
20'b01001111010110011101: color_data = 12'b111011101110;
20'b01001111010110011110: color_data = 12'b111011101110;
20'b01001111010110011111: color_data = 12'b111011101110;
20'b01001111010110100000: color_data = 12'b111011101110;
20'b01001111010110100001: color_data = 12'b111011101110;
20'b01001111010110100010: color_data = 12'b111011101110;
20'b01001111010110100011: color_data = 12'b111011101110;
20'b01001111010110100100: color_data = 12'b111011101110;
20'b01001111010110100101: color_data = 12'b111011101110;
20'b01001111010110100111: color_data = 12'b111011101110;
20'b01001111010110101000: color_data = 12'b111011101110;
20'b01001111010110101001: color_data = 12'b111011101110;
20'b01001111010110101010: color_data = 12'b111011101110;
20'b01001111010110101011: color_data = 12'b111011101110;
20'b01001111010110101100: color_data = 12'b111011101110;
20'b01001111010110101101: color_data = 12'b111011101110;
20'b01001111010110101110: color_data = 12'b111011101110;
20'b01001111010110101111: color_data = 12'b111011101110;
20'b01001111010110110000: color_data = 12'b111011101110;
20'b01001111010110111101: color_data = 12'b111011101110;
20'b01001111010110111110: color_data = 12'b111011101110;
20'b01001111010110111111: color_data = 12'b111011101110;
20'b01001111010111000000: color_data = 12'b111011101110;
20'b01001111010111000001: color_data = 12'b111011101110;
20'b01001111010111000010: color_data = 12'b111011101110;
20'b01001111010111000011: color_data = 12'b111011101110;
20'b01001111010111000100: color_data = 12'b111011101110;
20'b01001111010111000101: color_data = 12'b111011101110;
20'b01001111010111000110: color_data = 12'b111011101110;
20'b01001111010111001000: color_data = 12'b111011101110;
20'b01001111010111001001: color_data = 12'b111011101110;
20'b01001111010111001010: color_data = 12'b111011101110;
20'b01001111010111001011: color_data = 12'b111011101110;
20'b01001111010111001100: color_data = 12'b111011101110;
20'b01001111010111001101: color_data = 12'b111011101110;
20'b01001111010111001110: color_data = 12'b111011101110;
20'b01001111010111001111: color_data = 12'b111011101110;
20'b01001111010111010000: color_data = 12'b111011101110;
20'b01001111010111010001: color_data = 12'b111011101110;
20'b01001111100010010110: color_data = 12'b111011101110;
20'b01001111100010010111: color_data = 12'b111011101110;
20'b01001111100010011000: color_data = 12'b111011101110;
20'b01001111100010011001: color_data = 12'b111011101110;
20'b01001111100010011010: color_data = 12'b111011101110;
20'b01001111100010011011: color_data = 12'b111011101110;
20'b01001111100010011100: color_data = 12'b111011101110;
20'b01001111100010011101: color_data = 12'b111011101110;
20'b01001111100010011110: color_data = 12'b111011101110;
20'b01001111100010011111: color_data = 12'b111011101110;
20'b01001111100010100001: color_data = 12'b111011101110;
20'b01001111100010100010: color_data = 12'b111011101110;
20'b01001111100010100011: color_data = 12'b111011101110;
20'b01001111100010100100: color_data = 12'b111011101110;
20'b01001111100010100101: color_data = 12'b111011101110;
20'b01001111100010100110: color_data = 12'b111011101110;
20'b01001111100010100111: color_data = 12'b111011101110;
20'b01001111100010101000: color_data = 12'b111011101110;
20'b01001111100010101001: color_data = 12'b111011101110;
20'b01001111100010101010: color_data = 12'b111011101110;
20'b01001111100011001101: color_data = 12'b111011101110;
20'b01001111100011001110: color_data = 12'b111011101110;
20'b01001111100011001111: color_data = 12'b111011101110;
20'b01001111100011010000: color_data = 12'b111011101110;
20'b01001111100011010001: color_data = 12'b111011101110;
20'b01001111100011010010: color_data = 12'b111011101110;
20'b01001111100011010011: color_data = 12'b111011101110;
20'b01001111100011010100: color_data = 12'b111011101110;
20'b01001111100011010101: color_data = 12'b111011101110;
20'b01001111100011010110: color_data = 12'b111011101110;
20'b01001111100011011000: color_data = 12'b111011101110;
20'b01001111100011011001: color_data = 12'b111011101110;
20'b01001111100011011010: color_data = 12'b111011101110;
20'b01001111100011011011: color_data = 12'b111011101110;
20'b01001111100011011100: color_data = 12'b111011101110;
20'b01001111100011011101: color_data = 12'b111011101110;
20'b01001111100011011110: color_data = 12'b111011101110;
20'b01001111100011011111: color_data = 12'b111011101110;
20'b01001111100011100000: color_data = 12'b111011101110;
20'b01001111100011100001: color_data = 12'b111011101110;
20'b01001111100011101101: color_data = 12'b111011101110;
20'b01001111100011101110: color_data = 12'b111011101110;
20'b01001111100011101111: color_data = 12'b111011101110;
20'b01001111100011110000: color_data = 12'b111011101110;
20'b01001111100011110001: color_data = 12'b111011101110;
20'b01001111100011110010: color_data = 12'b111011101110;
20'b01001111100011110011: color_data = 12'b111011101110;
20'b01001111100011110100: color_data = 12'b111011101110;
20'b01001111100011110101: color_data = 12'b111011101110;
20'b01001111100011110110: color_data = 12'b111011101110;
20'b01001111100011111000: color_data = 12'b111011101110;
20'b01001111100011111001: color_data = 12'b111011101110;
20'b01001111100011111010: color_data = 12'b111011101110;
20'b01001111100011111011: color_data = 12'b111011101110;
20'b01001111100011111100: color_data = 12'b111011101110;
20'b01001111100011111101: color_data = 12'b111011101110;
20'b01001111100011111110: color_data = 12'b111011101110;
20'b01001111100011111111: color_data = 12'b111011101110;
20'b01001111100100000000: color_data = 12'b111011101110;
20'b01001111100100000001: color_data = 12'b111011101110;
20'b01001111100100000011: color_data = 12'b111011101110;
20'b01001111100100000100: color_data = 12'b111011101110;
20'b01001111100100000101: color_data = 12'b111011101110;
20'b01001111100100000110: color_data = 12'b111011101110;
20'b01001111100100000111: color_data = 12'b111011101110;
20'b01001111100100001000: color_data = 12'b111011101110;
20'b01001111100100001001: color_data = 12'b111011101110;
20'b01001111100100001010: color_data = 12'b111011101110;
20'b01001111100100001011: color_data = 12'b111011101110;
20'b01001111100100001100: color_data = 12'b111011101110;
20'b01001111100100011001: color_data = 12'b111011101110;
20'b01001111100100011010: color_data = 12'b111011101110;
20'b01001111100100011011: color_data = 12'b111011101110;
20'b01001111100100011100: color_data = 12'b111011101110;
20'b01001111100100011101: color_data = 12'b111011101110;
20'b01001111100100011110: color_data = 12'b111011101110;
20'b01001111100100011111: color_data = 12'b111011101110;
20'b01001111100100100000: color_data = 12'b111011101110;
20'b01001111100100100001: color_data = 12'b111011101110;
20'b01001111100100100010: color_data = 12'b111011101110;
20'b01001111100100100100: color_data = 12'b111011101110;
20'b01001111100100100101: color_data = 12'b111011101110;
20'b01001111100100100110: color_data = 12'b111011101110;
20'b01001111100100100111: color_data = 12'b111011101110;
20'b01001111100100101000: color_data = 12'b111011101110;
20'b01001111100100101001: color_data = 12'b111011101110;
20'b01001111100100101010: color_data = 12'b111011101110;
20'b01001111100100101011: color_data = 12'b111011101110;
20'b01001111100100101100: color_data = 12'b111011101110;
20'b01001111100100101101: color_data = 12'b111011101110;
20'b01001111100100101111: color_data = 12'b111011101110;
20'b01001111100100110000: color_data = 12'b111011101110;
20'b01001111100100110001: color_data = 12'b111011101110;
20'b01001111100100110010: color_data = 12'b111011101110;
20'b01001111100100110011: color_data = 12'b111011101110;
20'b01001111100100110100: color_data = 12'b111011101110;
20'b01001111100100110101: color_data = 12'b111011101110;
20'b01001111100100110110: color_data = 12'b111011101110;
20'b01001111100100110111: color_data = 12'b111011101110;
20'b01001111100100111000: color_data = 12'b111011101110;
20'b01001111100101000100: color_data = 12'b111011101110;
20'b01001111100101000101: color_data = 12'b111011101110;
20'b01001111100101000110: color_data = 12'b111011101110;
20'b01001111100101000111: color_data = 12'b111011101110;
20'b01001111100101001000: color_data = 12'b111011101110;
20'b01001111100101001001: color_data = 12'b111011101110;
20'b01001111100101001010: color_data = 12'b111011101110;
20'b01001111100101001011: color_data = 12'b111011101110;
20'b01001111100101001100: color_data = 12'b111011101110;
20'b01001111100101001101: color_data = 12'b111011101110;
20'b01001111100101001111: color_data = 12'b111011101110;
20'b01001111100101010000: color_data = 12'b111011101110;
20'b01001111100101010001: color_data = 12'b111011101110;
20'b01001111100101010010: color_data = 12'b111011101110;
20'b01001111100101010011: color_data = 12'b111011101110;
20'b01001111100101010100: color_data = 12'b111011101110;
20'b01001111100101010101: color_data = 12'b111011101110;
20'b01001111100101010110: color_data = 12'b111011101110;
20'b01001111100101010111: color_data = 12'b111011101110;
20'b01001111100101011000: color_data = 12'b111011101110;
20'b01001111100110011100: color_data = 12'b111011101110;
20'b01001111100110011101: color_data = 12'b111011101110;
20'b01001111100110011110: color_data = 12'b111011101110;
20'b01001111100110011111: color_data = 12'b111011101110;
20'b01001111100110100000: color_data = 12'b111011101110;
20'b01001111100110100001: color_data = 12'b111011101110;
20'b01001111100110100010: color_data = 12'b111011101110;
20'b01001111100110100011: color_data = 12'b111011101110;
20'b01001111100110100100: color_data = 12'b111011101110;
20'b01001111100110100101: color_data = 12'b111011101110;
20'b01001111100110100111: color_data = 12'b111011101110;
20'b01001111100110101000: color_data = 12'b111011101110;
20'b01001111100110101001: color_data = 12'b111011101110;
20'b01001111100110101010: color_data = 12'b111011101110;
20'b01001111100110101011: color_data = 12'b111011101110;
20'b01001111100110101100: color_data = 12'b111011101110;
20'b01001111100110101101: color_data = 12'b111011101110;
20'b01001111100110101110: color_data = 12'b111011101110;
20'b01001111100110101111: color_data = 12'b111011101110;
20'b01001111100110110000: color_data = 12'b111011101110;
20'b01001111100110111101: color_data = 12'b111011101110;
20'b01001111100110111110: color_data = 12'b111011101110;
20'b01001111100110111111: color_data = 12'b111011101110;
20'b01001111100111000000: color_data = 12'b111011101110;
20'b01001111100111000001: color_data = 12'b111011101110;
20'b01001111100111000010: color_data = 12'b111011101110;
20'b01001111100111000011: color_data = 12'b111011101110;
20'b01001111100111000100: color_data = 12'b111011101110;
20'b01001111100111000101: color_data = 12'b111011101110;
20'b01001111100111000110: color_data = 12'b111011101110;
20'b01001111100111001000: color_data = 12'b111011101110;
20'b01001111100111001001: color_data = 12'b111011101110;
20'b01001111100111001010: color_data = 12'b111011101110;
20'b01001111100111001011: color_data = 12'b111011101110;
20'b01001111100111001100: color_data = 12'b111011101110;
20'b01001111100111001101: color_data = 12'b111011101110;
20'b01001111100111001110: color_data = 12'b111011101110;
20'b01001111100111001111: color_data = 12'b111011101110;
20'b01001111100111010000: color_data = 12'b111011101110;
20'b01001111100111010001: color_data = 12'b111011101110;
20'b01001111110010010110: color_data = 12'b111011101110;
20'b01001111110010010111: color_data = 12'b111011101110;
20'b01001111110010011000: color_data = 12'b111011101110;
20'b01001111110010011001: color_data = 12'b111011101110;
20'b01001111110010011010: color_data = 12'b111011101110;
20'b01001111110010011011: color_data = 12'b111011101110;
20'b01001111110010011100: color_data = 12'b111011101110;
20'b01001111110010011101: color_data = 12'b111011101110;
20'b01001111110010011110: color_data = 12'b111011101110;
20'b01001111110010011111: color_data = 12'b111011101110;
20'b01001111110010100001: color_data = 12'b111011101110;
20'b01001111110010100010: color_data = 12'b111011101110;
20'b01001111110010100011: color_data = 12'b111011101110;
20'b01001111110010100100: color_data = 12'b111011101110;
20'b01001111110010100101: color_data = 12'b111011101110;
20'b01001111110010100110: color_data = 12'b111011101110;
20'b01001111110010100111: color_data = 12'b111011101110;
20'b01001111110010101000: color_data = 12'b111011101110;
20'b01001111110010101001: color_data = 12'b111011101110;
20'b01001111110010101010: color_data = 12'b111011101110;
20'b01001111110011001101: color_data = 12'b111011101110;
20'b01001111110011001110: color_data = 12'b111011101110;
20'b01001111110011001111: color_data = 12'b111011101110;
20'b01001111110011010000: color_data = 12'b111011101110;
20'b01001111110011010001: color_data = 12'b111011101110;
20'b01001111110011010010: color_data = 12'b111011101110;
20'b01001111110011010011: color_data = 12'b111011101110;
20'b01001111110011010100: color_data = 12'b111011101110;
20'b01001111110011010101: color_data = 12'b111011101110;
20'b01001111110011010110: color_data = 12'b111011101110;
20'b01001111110011011000: color_data = 12'b111011101110;
20'b01001111110011011001: color_data = 12'b111011101110;
20'b01001111110011011010: color_data = 12'b111011101110;
20'b01001111110011011011: color_data = 12'b111011101110;
20'b01001111110011011100: color_data = 12'b111011101110;
20'b01001111110011011101: color_data = 12'b111011101110;
20'b01001111110011011110: color_data = 12'b111011101110;
20'b01001111110011011111: color_data = 12'b111011101110;
20'b01001111110011100000: color_data = 12'b111011101110;
20'b01001111110011100001: color_data = 12'b111011101110;
20'b01001111110011101101: color_data = 12'b111011101110;
20'b01001111110011101110: color_data = 12'b111011101110;
20'b01001111110011101111: color_data = 12'b111011101110;
20'b01001111110011110000: color_data = 12'b111011101110;
20'b01001111110011110001: color_data = 12'b111011101110;
20'b01001111110011110010: color_data = 12'b111011101110;
20'b01001111110011110011: color_data = 12'b111011101110;
20'b01001111110011110100: color_data = 12'b111011101110;
20'b01001111110011110101: color_data = 12'b111011101110;
20'b01001111110011110110: color_data = 12'b111011101110;
20'b01001111110011111000: color_data = 12'b111011101110;
20'b01001111110011111001: color_data = 12'b111011101110;
20'b01001111110011111010: color_data = 12'b111011101110;
20'b01001111110011111011: color_data = 12'b111011101110;
20'b01001111110011111100: color_data = 12'b111011101110;
20'b01001111110011111101: color_data = 12'b111011101110;
20'b01001111110011111110: color_data = 12'b111011101110;
20'b01001111110011111111: color_data = 12'b111011101110;
20'b01001111110100000000: color_data = 12'b111011101110;
20'b01001111110100000001: color_data = 12'b111011101110;
20'b01001111110100000011: color_data = 12'b111011101110;
20'b01001111110100000100: color_data = 12'b111011101110;
20'b01001111110100000101: color_data = 12'b111011101110;
20'b01001111110100000110: color_data = 12'b111011101110;
20'b01001111110100000111: color_data = 12'b111011101110;
20'b01001111110100001000: color_data = 12'b111011101110;
20'b01001111110100001001: color_data = 12'b111011101110;
20'b01001111110100001010: color_data = 12'b111011101110;
20'b01001111110100001011: color_data = 12'b111011101110;
20'b01001111110100001100: color_data = 12'b111011101110;
20'b01001111110100011001: color_data = 12'b111011101110;
20'b01001111110100011010: color_data = 12'b111011101110;
20'b01001111110100011011: color_data = 12'b111011101110;
20'b01001111110100011100: color_data = 12'b111011101110;
20'b01001111110100011101: color_data = 12'b111011101110;
20'b01001111110100011110: color_data = 12'b111011101110;
20'b01001111110100011111: color_data = 12'b111011101110;
20'b01001111110100100000: color_data = 12'b111011101110;
20'b01001111110100100001: color_data = 12'b111011101110;
20'b01001111110100100010: color_data = 12'b111011101110;
20'b01001111110100100100: color_data = 12'b111011101110;
20'b01001111110100100101: color_data = 12'b111011101110;
20'b01001111110100100110: color_data = 12'b111011101110;
20'b01001111110100100111: color_data = 12'b111011101110;
20'b01001111110100101000: color_data = 12'b111011101110;
20'b01001111110100101001: color_data = 12'b111011101110;
20'b01001111110100101010: color_data = 12'b111011101110;
20'b01001111110100101011: color_data = 12'b111011101110;
20'b01001111110100101100: color_data = 12'b111011101110;
20'b01001111110100101101: color_data = 12'b111011101110;
20'b01001111110100101111: color_data = 12'b111011101110;
20'b01001111110100110000: color_data = 12'b111011101110;
20'b01001111110100110001: color_data = 12'b111011101110;
20'b01001111110100110010: color_data = 12'b111011101110;
20'b01001111110100110011: color_data = 12'b111011101110;
20'b01001111110100110100: color_data = 12'b111011101110;
20'b01001111110100110101: color_data = 12'b111011101110;
20'b01001111110100110110: color_data = 12'b111011101110;
20'b01001111110100110111: color_data = 12'b111011101110;
20'b01001111110100111000: color_data = 12'b111011101110;
20'b01001111110101000100: color_data = 12'b111011101110;
20'b01001111110101000101: color_data = 12'b111011101110;
20'b01001111110101000110: color_data = 12'b111011101110;
20'b01001111110101000111: color_data = 12'b111011101110;
20'b01001111110101001000: color_data = 12'b111011101110;
20'b01001111110101001001: color_data = 12'b111011101110;
20'b01001111110101001010: color_data = 12'b111011101110;
20'b01001111110101001011: color_data = 12'b111011101110;
20'b01001111110101001100: color_data = 12'b111011101110;
20'b01001111110101001101: color_data = 12'b111011101110;
20'b01001111110101001111: color_data = 12'b111011101110;
20'b01001111110101010000: color_data = 12'b111011101110;
20'b01001111110101010001: color_data = 12'b111011101110;
20'b01001111110101010010: color_data = 12'b111011101110;
20'b01001111110101010011: color_data = 12'b111011101110;
20'b01001111110101010100: color_data = 12'b111011101110;
20'b01001111110101010101: color_data = 12'b111011101110;
20'b01001111110101010110: color_data = 12'b111011101110;
20'b01001111110101010111: color_data = 12'b111011101110;
20'b01001111110101011000: color_data = 12'b111011101110;
20'b01001111110110011100: color_data = 12'b111011101110;
20'b01001111110110011101: color_data = 12'b111011101110;
20'b01001111110110011110: color_data = 12'b111011101110;
20'b01001111110110011111: color_data = 12'b111011101110;
20'b01001111110110100000: color_data = 12'b111011101110;
20'b01001111110110100001: color_data = 12'b111011101110;
20'b01001111110110100010: color_data = 12'b111011101110;
20'b01001111110110100011: color_data = 12'b111011101110;
20'b01001111110110100100: color_data = 12'b111011101110;
20'b01001111110110100101: color_data = 12'b111011101110;
20'b01001111110110100111: color_data = 12'b111011101110;
20'b01001111110110101000: color_data = 12'b111011101110;
20'b01001111110110101001: color_data = 12'b111011101110;
20'b01001111110110101010: color_data = 12'b111011101110;
20'b01001111110110101011: color_data = 12'b111011101110;
20'b01001111110110101100: color_data = 12'b111011101110;
20'b01001111110110101101: color_data = 12'b111011101110;
20'b01001111110110101110: color_data = 12'b111011101110;
20'b01001111110110101111: color_data = 12'b111011101110;
20'b01001111110110110000: color_data = 12'b111011101110;
20'b01001111110110111101: color_data = 12'b111011101110;
20'b01001111110110111110: color_data = 12'b111011101110;
20'b01001111110110111111: color_data = 12'b111011101110;
20'b01001111110111000000: color_data = 12'b111011101110;
20'b01001111110111000001: color_data = 12'b111011101110;
20'b01001111110111000010: color_data = 12'b111011101110;
20'b01001111110111000011: color_data = 12'b111011101110;
20'b01001111110111000100: color_data = 12'b111011101110;
20'b01001111110111000101: color_data = 12'b111011101110;
20'b01001111110111000110: color_data = 12'b111011101110;
20'b01001111110111001000: color_data = 12'b111011101110;
20'b01001111110111001001: color_data = 12'b111011101110;
20'b01001111110111001010: color_data = 12'b111011101110;
20'b01001111110111001011: color_data = 12'b111011101110;
20'b01001111110111001100: color_data = 12'b111011101110;
20'b01001111110111001101: color_data = 12'b111011101110;
20'b01001111110111001110: color_data = 12'b111011101110;
20'b01001111110111001111: color_data = 12'b111011101110;
20'b01001111110111010000: color_data = 12'b111011101110;
20'b01001111110111010001: color_data = 12'b111011101110;
20'b01010000000010010110: color_data = 12'b111011101110;
20'b01010000000010010111: color_data = 12'b111011101110;
20'b01010000000010011000: color_data = 12'b111011101110;
20'b01010000000010011001: color_data = 12'b111011101110;
20'b01010000000010011010: color_data = 12'b111011101110;
20'b01010000000010011011: color_data = 12'b111011101110;
20'b01010000000010011100: color_data = 12'b111011101110;
20'b01010000000010011101: color_data = 12'b111011101110;
20'b01010000000010011110: color_data = 12'b111011101110;
20'b01010000000010011111: color_data = 12'b111011101110;
20'b01010000000010100001: color_data = 12'b111011101110;
20'b01010000000010100010: color_data = 12'b111011101110;
20'b01010000000010100011: color_data = 12'b111011101110;
20'b01010000000010100100: color_data = 12'b111011101110;
20'b01010000000010100101: color_data = 12'b111011101110;
20'b01010000000010100110: color_data = 12'b111011101110;
20'b01010000000010100111: color_data = 12'b111011101110;
20'b01010000000010101000: color_data = 12'b111011101110;
20'b01010000000010101001: color_data = 12'b111011101110;
20'b01010000000010101010: color_data = 12'b111011101110;
20'b01010000000011001101: color_data = 12'b111011101110;
20'b01010000000011001110: color_data = 12'b111011101110;
20'b01010000000011001111: color_data = 12'b111011101110;
20'b01010000000011010000: color_data = 12'b111011101110;
20'b01010000000011010001: color_data = 12'b111011101110;
20'b01010000000011010010: color_data = 12'b111011101110;
20'b01010000000011010011: color_data = 12'b111011101110;
20'b01010000000011010100: color_data = 12'b111011101110;
20'b01010000000011010101: color_data = 12'b111011101110;
20'b01010000000011010110: color_data = 12'b111011101110;
20'b01010000000011011000: color_data = 12'b111011101110;
20'b01010000000011011001: color_data = 12'b111011101110;
20'b01010000000011011010: color_data = 12'b111011101110;
20'b01010000000011011011: color_data = 12'b111011101110;
20'b01010000000011011100: color_data = 12'b111011101110;
20'b01010000000011011101: color_data = 12'b111011101110;
20'b01010000000011011110: color_data = 12'b111011101110;
20'b01010000000011011111: color_data = 12'b111011101110;
20'b01010000000011100000: color_data = 12'b111011101110;
20'b01010000000011100001: color_data = 12'b111011101110;
20'b01010000000011101101: color_data = 12'b111011101110;
20'b01010000000011101110: color_data = 12'b111011101110;
20'b01010000000011101111: color_data = 12'b111011101110;
20'b01010000000011110000: color_data = 12'b111011101110;
20'b01010000000011110001: color_data = 12'b111011101110;
20'b01010000000011110010: color_data = 12'b111011101110;
20'b01010000000011110011: color_data = 12'b111011101110;
20'b01010000000011110100: color_data = 12'b111011101110;
20'b01010000000011110101: color_data = 12'b111011101110;
20'b01010000000011110110: color_data = 12'b111011101110;
20'b01010000000011111000: color_data = 12'b111011101110;
20'b01010000000011111001: color_data = 12'b111011101110;
20'b01010000000011111010: color_data = 12'b111011101110;
20'b01010000000011111011: color_data = 12'b111011101110;
20'b01010000000011111100: color_data = 12'b111011101110;
20'b01010000000011111101: color_data = 12'b111011101110;
20'b01010000000011111110: color_data = 12'b111011101110;
20'b01010000000011111111: color_data = 12'b111011101110;
20'b01010000000100000000: color_data = 12'b111011101110;
20'b01010000000100000001: color_data = 12'b111011101110;
20'b01010000000100000011: color_data = 12'b111011101110;
20'b01010000000100000100: color_data = 12'b111011101110;
20'b01010000000100000101: color_data = 12'b111011101110;
20'b01010000000100000110: color_data = 12'b111011101110;
20'b01010000000100000111: color_data = 12'b111011101110;
20'b01010000000100001000: color_data = 12'b111011101110;
20'b01010000000100001001: color_data = 12'b111011101110;
20'b01010000000100001010: color_data = 12'b111011101110;
20'b01010000000100001011: color_data = 12'b111011101110;
20'b01010000000100001100: color_data = 12'b111011101110;
20'b01010000000100011001: color_data = 12'b111011101110;
20'b01010000000100011010: color_data = 12'b111011101110;
20'b01010000000100011011: color_data = 12'b111011101110;
20'b01010000000100011100: color_data = 12'b111011101110;
20'b01010000000100011101: color_data = 12'b111011101110;
20'b01010000000100011110: color_data = 12'b111011101110;
20'b01010000000100011111: color_data = 12'b111011101110;
20'b01010000000100100000: color_data = 12'b111011101110;
20'b01010000000100100001: color_data = 12'b111011101110;
20'b01010000000100100010: color_data = 12'b111011101110;
20'b01010000000100100100: color_data = 12'b111011101110;
20'b01010000000100100101: color_data = 12'b111011101110;
20'b01010000000100100110: color_data = 12'b111011101110;
20'b01010000000100100111: color_data = 12'b111011101110;
20'b01010000000100101000: color_data = 12'b111011101110;
20'b01010000000100101001: color_data = 12'b111011101110;
20'b01010000000100101010: color_data = 12'b111011101110;
20'b01010000000100101011: color_data = 12'b111011101110;
20'b01010000000100101100: color_data = 12'b111011101110;
20'b01010000000100101101: color_data = 12'b111011101110;
20'b01010000000100101111: color_data = 12'b111011101110;
20'b01010000000100110000: color_data = 12'b111011101110;
20'b01010000000100110001: color_data = 12'b111011101110;
20'b01010000000100110010: color_data = 12'b111011101110;
20'b01010000000100110011: color_data = 12'b111011101110;
20'b01010000000100110100: color_data = 12'b111011101110;
20'b01010000000100110101: color_data = 12'b111011101110;
20'b01010000000100110110: color_data = 12'b111011101110;
20'b01010000000100110111: color_data = 12'b111011101110;
20'b01010000000100111000: color_data = 12'b111011101110;
20'b01010000000101000100: color_data = 12'b111011101110;
20'b01010000000101000101: color_data = 12'b111011101110;
20'b01010000000101000110: color_data = 12'b111011101110;
20'b01010000000101000111: color_data = 12'b111011101110;
20'b01010000000101001000: color_data = 12'b111011101110;
20'b01010000000101001001: color_data = 12'b111011101110;
20'b01010000000101001010: color_data = 12'b111011101110;
20'b01010000000101001011: color_data = 12'b111011101110;
20'b01010000000101001100: color_data = 12'b111011101110;
20'b01010000000101001101: color_data = 12'b111011101110;
20'b01010000000101001111: color_data = 12'b111011101110;
20'b01010000000101010000: color_data = 12'b111011101110;
20'b01010000000101010001: color_data = 12'b111011101110;
20'b01010000000101010010: color_data = 12'b111011101110;
20'b01010000000101010011: color_data = 12'b111011101110;
20'b01010000000101010100: color_data = 12'b111011101110;
20'b01010000000101010101: color_data = 12'b111011101110;
20'b01010000000101010110: color_data = 12'b111011101110;
20'b01010000000101010111: color_data = 12'b111011101110;
20'b01010000000101011000: color_data = 12'b111011101110;
20'b01010000000110011100: color_data = 12'b111011101110;
20'b01010000000110011101: color_data = 12'b111011101110;
20'b01010000000110011110: color_data = 12'b111011101110;
20'b01010000000110011111: color_data = 12'b111011101110;
20'b01010000000110100000: color_data = 12'b111011101110;
20'b01010000000110100001: color_data = 12'b111011101110;
20'b01010000000110100010: color_data = 12'b111011101110;
20'b01010000000110100011: color_data = 12'b111011101110;
20'b01010000000110100100: color_data = 12'b111011101110;
20'b01010000000110100101: color_data = 12'b111011101110;
20'b01010000000110100111: color_data = 12'b111011101110;
20'b01010000000110101000: color_data = 12'b111011101110;
20'b01010000000110101001: color_data = 12'b111011101110;
20'b01010000000110101010: color_data = 12'b111011101110;
20'b01010000000110101011: color_data = 12'b111011101110;
20'b01010000000110101100: color_data = 12'b111011101110;
20'b01010000000110101101: color_data = 12'b111011101110;
20'b01010000000110101110: color_data = 12'b111011101110;
20'b01010000000110101111: color_data = 12'b111011101110;
20'b01010000000110110000: color_data = 12'b111011101110;
20'b01010000000110111101: color_data = 12'b111011101110;
20'b01010000000110111110: color_data = 12'b111011101110;
20'b01010000000110111111: color_data = 12'b111011101110;
20'b01010000000111000000: color_data = 12'b111011101110;
20'b01010000000111000001: color_data = 12'b111011101110;
20'b01010000000111000010: color_data = 12'b111011101110;
20'b01010000000111000011: color_data = 12'b111011101110;
20'b01010000000111000100: color_data = 12'b111011101110;
20'b01010000000111000101: color_data = 12'b111011101110;
20'b01010000000111000110: color_data = 12'b111011101110;
20'b01010000000111001000: color_data = 12'b111011101110;
20'b01010000000111001001: color_data = 12'b111011101110;
20'b01010000000111001010: color_data = 12'b111011101110;
20'b01010000000111001011: color_data = 12'b111011101110;
20'b01010000000111001100: color_data = 12'b111011101110;
20'b01010000000111001101: color_data = 12'b111011101110;
20'b01010000000111001110: color_data = 12'b111011101110;
20'b01010000000111001111: color_data = 12'b111011101110;
20'b01010000000111010000: color_data = 12'b111011101110;
20'b01010000000111010001: color_data = 12'b111011101110;
20'b01010000100010100001: color_data = 12'b111011101110;
20'b01010000100010100010: color_data = 12'b111011101110;
20'b01010000100010100011: color_data = 12'b111011101110;
20'b01010000100010100100: color_data = 12'b111011101110;
20'b01010000100010100101: color_data = 12'b111011101110;
20'b01010000100010100110: color_data = 12'b111011101110;
20'b01010000100010100111: color_data = 12'b111011101110;
20'b01010000100010101000: color_data = 12'b111011101110;
20'b01010000100010101001: color_data = 12'b111011101110;
20'b01010000100010101010: color_data = 12'b111011101110;
20'b01010000100010101100: color_data = 12'b111011101110;
20'b01010000100010101101: color_data = 12'b111011101110;
20'b01010000100010101110: color_data = 12'b111011101110;
20'b01010000100010101111: color_data = 12'b111011101110;
20'b01010000100010110000: color_data = 12'b111011101110;
20'b01010000100010110001: color_data = 12'b111011101110;
20'b01010000100010110010: color_data = 12'b111011101110;
20'b01010000100010110011: color_data = 12'b111011101110;
20'b01010000100010110100: color_data = 12'b111011101110;
20'b01010000100010110101: color_data = 12'b111011101110;
20'b01010000100010110111: color_data = 12'b111011101110;
20'b01010000100010111000: color_data = 12'b111011101110;
20'b01010000100010111001: color_data = 12'b111011101110;
20'b01010000100010111010: color_data = 12'b111011101110;
20'b01010000100010111011: color_data = 12'b111011101110;
20'b01010000100010111100: color_data = 12'b111011101110;
20'b01010000100010111101: color_data = 12'b111011101110;
20'b01010000100010111110: color_data = 12'b111011101110;
20'b01010000100010111111: color_data = 12'b111011101110;
20'b01010000100011000000: color_data = 12'b111011101110;
20'b01010000100011000010: color_data = 12'b111011101110;
20'b01010000100011000011: color_data = 12'b111011101110;
20'b01010000100011000100: color_data = 12'b111011101110;
20'b01010000100011000101: color_data = 12'b111011101110;
20'b01010000100011000110: color_data = 12'b111011101110;
20'b01010000100011000111: color_data = 12'b111011101110;
20'b01010000100011001000: color_data = 12'b111011101110;
20'b01010000100011001001: color_data = 12'b111011101110;
20'b01010000100011001010: color_data = 12'b111011101110;
20'b01010000100011001011: color_data = 12'b111011101110;
20'b01010000100011001101: color_data = 12'b111011101110;
20'b01010000100011001110: color_data = 12'b111011101110;
20'b01010000100011001111: color_data = 12'b111011101110;
20'b01010000100011010000: color_data = 12'b111011101110;
20'b01010000100011010001: color_data = 12'b111011101110;
20'b01010000100011010010: color_data = 12'b111011101110;
20'b01010000100011010011: color_data = 12'b111011101110;
20'b01010000100011010100: color_data = 12'b111011101110;
20'b01010000100011010101: color_data = 12'b111011101110;
20'b01010000100011010110: color_data = 12'b111011101110;
20'b01010000100011111000: color_data = 12'b111011101110;
20'b01010000100011111001: color_data = 12'b111011101110;
20'b01010000100011111010: color_data = 12'b111011101110;
20'b01010000100011111011: color_data = 12'b111011101110;
20'b01010000100011111100: color_data = 12'b111011101110;
20'b01010000100011111101: color_data = 12'b111011101110;
20'b01010000100011111110: color_data = 12'b111011101110;
20'b01010000100011111111: color_data = 12'b111011101110;
20'b01010000100100000000: color_data = 12'b111011101110;
20'b01010000100100000001: color_data = 12'b111011101110;
20'b01010000100100000011: color_data = 12'b111011101110;
20'b01010000100100000100: color_data = 12'b111011101110;
20'b01010000100100000101: color_data = 12'b111011101110;
20'b01010000100100000110: color_data = 12'b111011101110;
20'b01010000100100000111: color_data = 12'b111011101110;
20'b01010000100100001000: color_data = 12'b111011101110;
20'b01010000100100001001: color_data = 12'b111011101110;
20'b01010000100100001010: color_data = 12'b111011101110;
20'b01010000100100001011: color_data = 12'b111011101110;
20'b01010000100100001100: color_data = 12'b111011101110;
20'b01010000100100001110: color_data = 12'b111011101110;
20'b01010000100100001111: color_data = 12'b111011101110;
20'b01010000100100010000: color_data = 12'b111011101110;
20'b01010000100100010001: color_data = 12'b111011101110;
20'b01010000100100010010: color_data = 12'b111011101110;
20'b01010000100100010011: color_data = 12'b111011101110;
20'b01010000100100010100: color_data = 12'b111011101110;
20'b01010000100100010101: color_data = 12'b111011101110;
20'b01010000100100010110: color_data = 12'b111011101110;
20'b01010000100100010111: color_data = 12'b111011101110;
20'b01010000100100011001: color_data = 12'b111011101110;
20'b01010000100100011010: color_data = 12'b111011101110;
20'b01010000100100011011: color_data = 12'b111011101110;
20'b01010000100100011100: color_data = 12'b111011101110;
20'b01010000100100011101: color_data = 12'b111011101110;
20'b01010000100100011110: color_data = 12'b111011101110;
20'b01010000100100011111: color_data = 12'b111011101110;
20'b01010000100100100000: color_data = 12'b111011101110;
20'b01010000100100100001: color_data = 12'b111011101110;
20'b01010000100100100010: color_data = 12'b111011101110;
20'b01010000100100100100: color_data = 12'b111011101110;
20'b01010000100100100101: color_data = 12'b111011101110;
20'b01010000100100100110: color_data = 12'b111011101110;
20'b01010000100100100111: color_data = 12'b111011101110;
20'b01010000100100101000: color_data = 12'b111011101110;
20'b01010000100100101001: color_data = 12'b111011101110;
20'b01010000100100101010: color_data = 12'b111011101110;
20'b01010000100100101011: color_data = 12'b111011101110;
20'b01010000100100101100: color_data = 12'b111011101110;
20'b01010000100100101101: color_data = 12'b111011101110;
20'b01010000100101000100: color_data = 12'b111011101110;
20'b01010000100101000101: color_data = 12'b111011101110;
20'b01010000100101000110: color_data = 12'b111011101110;
20'b01010000100101000111: color_data = 12'b111011101110;
20'b01010000100101001000: color_data = 12'b111011101110;
20'b01010000100101001001: color_data = 12'b111011101110;
20'b01010000100101001010: color_data = 12'b111011101110;
20'b01010000100101001011: color_data = 12'b111011101110;
20'b01010000100101001100: color_data = 12'b111011101110;
20'b01010000100101001101: color_data = 12'b111011101110;
20'b01010000100101001111: color_data = 12'b111011101110;
20'b01010000100101010000: color_data = 12'b111011101110;
20'b01010000100101010001: color_data = 12'b111011101110;
20'b01010000100101010010: color_data = 12'b111011101110;
20'b01010000100101010011: color_data = 12'b111011101110;
20'b01010000100101010100: color_data = 12'b111011101110;
20'b01010000100101010101: color_data = 12'b111011101110;
20'b01010000100101010110: color_data = 12'b111011101110;
20'b01010000100101010111: color_data = 12'b111011101110;
20'b01010000100101011000: color_data = 12'b111011101110;
20'b01010000100101011010: color_data = 12'b111011101110;
20'b01010000100101011011: color_data = 12'b111011101110;
20'b01010000100101011100: color_data = 12'b111011101110;
20'b01010000100101011101: color_data = 12'b111011101110;
20'b01010000100101011110: color_data = 12'b111011101110;
20'b01010000100101011111: color_data = 12'b111011101110;
20'b01010000100101100000: color_data = 12'b111011101110;
20'b01010000100101100001: color_data = 12'b111011101110;
20'b01010000100101100010: color_data = 12'b111011101110;
20'b01010000100101100011: color_data = 12'b111011101110;
20'b01010000100101100101: color_data = 12'b111011101110;
20'b01010000100101100110: color_data = 12'b111011101110;
20'b01010000100101100111: color_data = 12'b111011101110;
20'b01010000100101101000: color_data = 12'b111011101110;
20'b01010000100101101001: color_data = 12'b111011101110;
20'b01010000100101101010: color_data = 12'b111011101110;
20'b01010000100101101011: color_data = 12'b111011101110;
20'b01010000100101101100: color_data = 12'b111011101110;
20'b01010000100101101101: color_data = 12'b111011101110;
20'b01010000100101101110: color_data = 12'b111011101110;
20'b01010000100101110000: color_data = 12'b111011101110;
20'b01010000100101110001: color_data = 12'b111011101110;
20'b01010000100101110010: color_data = 12'b111011101110;
20'b01010000100101110011: color_data = 12'b111011101110;
20'b01010000100101110100: color_data = 12'b111011101110;
20'b01010000100101110101: color_data = 12'b111011101110;
20'b01010000100101110110: color_data = 12'b111011101110;
20'b01010000100101110111: color_data = 12'b111011101110;
20'b01010000100101111000: color_data = 12'b111011101110;
20'b01010000100101111001: color_data = 12'b111011101110;
20'b01010000100101111011: color_data = 12'b111011101110;
20'b01010000100101111100: color_data = 12'b111011101110;
20'b01010000100101111101: color_data = 12'b111011101110;
20'b01010000100101111110: color_data = 12'b111011101110;
20'b01010000100101111111: color_data = 12'b111011101110;
20'b01010000100110000000: color_data = 12'b111011101110;
20'b01010000100110000001: color_data = 12'b111011101110;
20'b01010000100110000010: color_data = 12'b111011101110;
20'b01010000100110000011: color_data = 12'b111011101110;
20'b01010000100110000100: color_data = 12'b111011101110;
20'b01010000100110000110: color_data = 12'b111011101110;
20'b01010000100110000111: color_data = 12'b111011101110;
20'b01010000100110001000: color_data = 12'b111011101110;
20'b01010000100110001001: color_data = 12'b111011101110;
20'b01010000100110001010: color_data = 12'b111011101110;
20'b01010000100110001011: color_data = 12'b111011101110;
20'b01010000100110001100: color_data = 12'b111011101110;
20'b01010000100110001101: color_data = 12'b111011101110;
20'b01010000100110001110: color_data = 12'b111011101110;
20'b01010000100110001111: color_data = 12'b111011101110;
20'b01010000100110011100: color_data = 12'b111011101110;
20'b01010000100110011101: color_data = 12'b111011101110;
20'b01010000100110011110: color_data = 12'b111011101110;
20'b01010000100110011111: color_data = 12'b111011101110;
20'b01010000100110100000: color_data = 12'b111011101110;
20'b01010000100110100001: color_data = 12'b111011101110;
20'b01010000100110100010: color_data = 12'b111011101110;
20'b01010000100110100011: color_data = 12'b111011101110;
20'b01010000100110100100: color_data = 12'b111011101110;
20'b01010000100110100101: color_data = 12'b111011101110;
20'b01010000100110100111: color_data = 12'b111011101110;
20'b01010000100110101000: color_data = 12'b111011101110;
20'b01010000100110101001: color_data = 12'b111011101110;
20'b01010000100110101010: color_data = 12'b111011101110;
20'b01010000100110101011: color_data = 12'b111011101110;
20'b01010000100110101100: color_data = 12'b111011101110;
20'b01010000100110101101: color_data = 12'b111011101110;
20'b01010000100110101110: color_data = 12'b111011101110;
20'b01010000100110101111: color_data = 12'b111011101110;
20'b01010000100110110000: color_data = 12'b111011101110;
20'b01010000100111001000: color_data = 12'b111011101110;
20'b01010000100111001001: color_data = 12'b111011101110;
20'b01010000100111001010: color_data = 12'b111011101110;
20'b01010000100111001011: color_data = 12'b111011101110;
20'b01010000100111001100: color_data = 12'b111011101110;
20'b01010000100111001101: color_data = 12'b111011101110;
20'b01010000100111001110: color_data = 12'b111011101110;
20'b01010000100111001111: color_data = 12'b111011101110;
20'b01010000100111010000: color_data = 12'b111011101110;
20'b01010000100111010001: color_data = 12'b111011101110;
20'b01010000100111010011: color_data = 12'b111011101110;
20'b01010000100111010100: color_data = 12'b111011101110;
20'b01010000100111010101: color_data = 12'b111011101110;
20'b01010000100111010110: color_data = 12'b111011101110;
20'b01010000100111010111: color_data = 12'b111011101110;
20'b01010000100111011000: color_data = 12'b111011101110;
20'b01010000100111011001: color_data = 12'b111011101110;
20'b01010000100111011010: color_data = 12'b111011101110;
20'b01010000100111011011: color_data = 12'b111011101110;
20'b01010000100111011100: color_data = 12'b111011101110;
20'b01010000110010100001: color_data = 12'b111011101110;
20'b01010000110010100010: color_data = 12'b111011101110;
20'b01010000110010100011: color_data = 12'b111011101110;
20'b01010000110010100100: color_data = 12'b111011101110;
20'b01010000110010100101: color_data = 12'b111011101110;
20'b01010000110010100110: color_data = 12'b111011101110;
20'b01010000110010100111: color_data = 12'b111011101110;
20'b01010000110010101000: color_data = 12'b111011101110;
20'b01010000110010101001: color_data = 12'b111011101110;
20'b01010000110010101010: color_data = 12'b111011101110;
20'b01010000110010101100: color_data = 12'b111011101110;
20'b01010000110010101101: color_data = 12'b111011101110;
20'b01010000110010101110: color_data = 12'b111011101110;
20'b01010000110010101111: color_data = 12'b111011101110;
20'b01010000110010110000: color_data = 12'b111011101110;
20'b01010000110010110001: color_data = 12'b111011101110;
20'b01010000110010110010: color_data = 12'b111011101110;
20'b01010000110010110011: color_data = 12'b111011101110;
20'b01010000110010110100: color_data = 12'b111011101110;
20'b01010000110010110101: color_data = 12'b111011101110;
20'b01010000110010110111: color_data = 12'b111011101110;
20'b01010000110010111000: color_data = 12'b111011101110;
20'b01010000110010111001: color_data = 12'b111011101110;
20'b01010000110010111010: color_data = 12'b111011101110;
20'b01010000110010111011: color_data = 12'b111011101110;
20'b01010000110010111100: color_data = 12'b111011101110;
20'b01010000110010111101: color_data = 12'b111011101110;
20'b01010000110010111110: color_data = 12'b111011101110;
20'b01010000110010111111: color_data = 12'b111011101110;
20'b01010000110011000000: color_data = 12'b111011101110;
20'b01010000110011000010: color_data = 12'b111011101110;
20'b01010000110011000011: color_data = 12'b111011101110;
20'b01010000110011000100: color_data = 12'b111011101110;
20'b01010000110011000101: color_data = 12'b111011101110;
20'b01010000110011000110: color_data = 12'b111011101110;
20'b01010000110011000111: color_data = 12'b111011101110;
20'b01010000110011001000: color_data = 12'b111011101110;
20'b01010000110011001001: color_data = 12'b111011101110;
20'b01010000110011001010: color_data = 12'b111011101110;
20'b01010000110011001011: color_data = 12'b111011101110;
20'b01010000110011001101: color_data = 12'b111011101110;
20'b01010000110011001110: color_data = 12'b111011101110;
20'b01010000110011001111: color_data = 12'b111011101110;
20'b01010000110011010000: color_data = 12'b111011101110;
20'b01010000110011010001: color_data = 12'b111011101110;
20'b01010000110011010010: color_data = 12'b111011101110;
20'b01010000110011010011: color_data = 12'b111011101110;
20'b01010000110011010100: color_data = 12'b111011101110;
20'b01010000110011010101: color_data = 12'b111011101110;
20'b01010000110011010110: color_data = 12'b111011101110;
20'b01010000110011111000: color_data = 12'b111011101110;
20'b01010000110011111001: color_data = 12'b111011101110;
20'b01010000110011111010: color_data = 12'b111011101110;
20'b01010000110011111011: color_data = 12'b111011101110;
20'b01010000110011111100: color_data = 12'b111011101110;
20'b01010000110011111101: color_data = 12'b111011101110;
20'b01010000110011111110: color_data = 12'b111011101110;
20'b01010000110011111111: color_data = 12'b111011101110;
20'b01010000110100000000: color_data = 12'b111011101110;
20'b01010000110100000001: color_data = 12'b111011101110;
20'b01010000110100000011: color_data = 12'b111011101110;
20'b01010000110100000100: color_data = 12'b111011101110;
20'b01010000110100000101: color_data = 12'b111011101110;
20'b01010000110100000110: color_data = 12'b111011101110;
20'b01010000110100000111: color_data = 12'b111011101110;
20'b01010000110100001000: color_data = 12'b111011101110;
20'b01010000110100001001: color_data = 12'b111011101110;
20'b01010000110100001010: color_data = 12'b111011101110;
20'b01010000110100001011: color_data = 12'b111011101110;
20'b01010000110100001100: color_data = 12'b111011101110;
20'b01010000110100001110: color_data = 12'b111011101110;
20'b01010000110100001111: color_data = 12'b111011101110;
20'b01010000110100010000: color_data = 12'b111011101110;
20'b01010000110100010001: color_data = 12'b111011101110;
20'b01010000110100010010: color_data = 12'b111011101110;
20'b01010000110100010011: color_data = 12'b111011101110;
20'b01010000110100010100: color_data = 12'b111011101110;
20'b01010000110100010101: color_data = 12'b111011101110;
20'b01010000110100010110: color_data = 12'b111011101110;
20'b01010000110100010111: color_data = 12'b111011101110;
20'b01010000110100011001: color_data = 12'b111011101110;
20'b01010000110100011010: color_data = 12'b111011101110;
20'b01010000110100011011: color_data = 12'b111011101110;
20'b01010000110100011100: color_data = 12'b111011101110;
20'b01010000110100011101: color_data = 12'b111011101110;
20'b01010000110100011110: color_data = 12'b111011101110;
20'b01010000110100011111: color_data = 12'b111011101110;
20'b01010000110100100000: color_data = 12'b111011101110;
20'b01010000110100100001: color_data = 12'b111011101110;
20'b01010000110100100010: color_data = 12'b111011101110;
20'b01010000110100100100: color_data = 12'b111011101110;
20'b01010000110100100101: color_data = 12'b111011101110;
20'b01010000110100100110: color_data = 12'b111011101110;
20'b01010000110100100111: color_data = 12'b111011101110;
20'b01010000110100101000: color_data = 12'b111011101110;
20'b01010000110100101001: color_data = 12'b111011101110;
20'b01010000110100101010: color_data = 12'b111011101110;
20'b01010000110100101011: color_data = 12'b111011101110;
20'b01010000110100101100: color_data = 12'b111011101110;
20'b01010000110100101101: color_data = 12'b111011101110;
20'b01010000110101000100: color_data = 12'b111011101110;
20'b01010000110101000101: color_data = 12'b111011101110;
20'b01010000110101000110: color_data = 12'b111011101110;
20'b01010000110101000111: color_data = 12'b111011101110;
20'b01010000110101001000: color_data = 12'b111011101110;
20'b01010000110101001001: color_data = 12'b111011101110;
20'b01010000110101001010: color_data = 12'b111011101110;
20'b01010000110101001011: color_data = 12'b111011101110;
20'b01010000110101001100: color_data = 12'b111011101110;
20'b01010000110101001101: color_data = 12'b111011101110;
20'b01010000110101001111: color_data = 12'b111011101110;
20'b01010000110101010000: color_data = 12'b111011101110;
20'b01010000110101010001: color_data = 12'b111011101110;
20'b01010000110101010010: color_data = 12'b111011101110;
20'b01010000110101010011: color_data = 12'b111011101110;
20'b01010000110101010100: color_data = 12'b111011101110;
20'b01010000110101010101: color_data = 12'b111011101110;
20'b01010000110101010110: color_data = 12'b111011101110;
20'b01010000110101010111: color_data = 12'b111011101110;
20'b01010000110101011000: color_data = 12'b111011101110;
20'b01010000110101011010: color_data = 12'b111011101110;
20'b01010000110101011011: color_data = 12'b111011101110;
20'b01010000110101011100: color_data = 12'b111011101110;
20'b01010000110101011101: color_data = 12'b111011101110;
20'b01010000110101011110: color_data = 12'b111011101110;
20'b01010000110101011111: color_data = 12'b111011101110;
20'b01010000110101100000: color_data = 12'b111011101110;
20'b01010000110101100001: color_data = 12'b111011101110;
20'b01010000110101100010: color_data = 12'b111011101110;
20'b01010000110101100011: color_data = 12'b111011101110;
20'b01010000110101100101: color_data = 12'b111011101110;
20'b01010000110101100110: color_data = 12'b111011101110;
20'b01010000110101100111: color_data = 12'b111011101110;
20'b01010000110101101000: color_data = 12'b111011101110;
20'b01010000110101101001: color_data = 12'b111011101110;
20'b01010000110101101010: color_data = 12'b111011101110;
20'b01010000110101101011: color_data = 12'b111011101110;
20'b01010000110101101100: color_data = 12'b111011101110;
20'b01010000110101101101: color_data = 12'b111011101110;
20'b01010000110101101110: color_data = 12'b111011101110;
20'b01010000110101110000: color_data = 12'b111011101110;
20'b01010000110101110001: color_data = 12'b111011101110;
20'b01010000110101110010: color_data = 12'b111011101110;
20'b01010000110101110011: color_data = 12'b111011101110;
20'b01010000110101110100: color_data = 12'b111011101110;
20'b01010000110101110101: color_data = 12'b111011101110;
20'b01010000110101110110: color_data = 12'b111011101110;
20'b01010000110101110111: color_data = 12'b111011101110;
20'b01010000110101111000: color_data = 12'b111011101110;
20'b01010000110101111001: color_data = 12'b111011101110;
20'b01010000110101111011: color_data = 12'b111011101110;
20'b01010000110101111100: color_data = 12'b111011101110;
20'b01010000110101111101: color_data = 12'b111011101110;
20'b01010000110101111110: color_data = 12'b111011101110;
20'b01010000110101111111: color_data = 12'b111011101110;
20'b01010000110110000000: color_data = 12'b111011101110;
20'b01010000110110000001: color_data = 12'b111011101110;
20'b01010000110110000010: color_data = 12'b111011101110;
20'b01010000110110000011: color_data = 12'b111011101110;
20'b01010000110110000100: color_data = 12'b111011101110;
20'b01010000110110000110: color_data = 12'b111011101110;
20'b01010000110110000111: color_data = 12'b111011101110;
20'b01010000110110001000: color_data = 12'b111011101110;
20'b01010000110110001001: color_data = 12'b111011101110;
20'b01010000110110001010: color_data = 12'b111011101110;
20'b01010000110110001011: color_data = 12'b111011101110;
20'b01010000110110001100: color_data = 12'b111011101110;
20'b01010000110110001101: color_data = 12'b111011101110;
20'b01010000110110001110: color_data = 12'b111011101110;
20'b01010000110110001111: color_data = 12'b111011101110;
20'b01010000110110011100: color_data = 12'b111011101110;
20'b01010000110110011101: color_data = 12'b111011101110;
20'b01010000110110011110: color_data = 12'b111011101110;
20'b01010000110110011111: color_data = 12'b111011101110;
20'b01010000110110100000: color_data = 12'b111011101110;
20'b01010000110110100001: color_data = 12'b111011101110;
20'b01010000110110100010: color_data = 12'b111011101110;
20'b01010000110110100011: color_data = 12'b111011101110;
20'b01010000110110100100: color_data = 12'b111011101110;
20'b01010000110110100101: color_data = 12'b111011101110;
20'b01010000110110100111: color_data = 12'b111011101110;
20'b01010000110110101000: color_data = 12'b111011101110;
20'b01010000110110101001: color_data = 12'b111011101110;
20'b01010000110110101010: color_data = 12'b111011101110;
20'b01010000110110101011: color_data = 12'b111011101110;
20'b01010000110110101100: color_data = 12'b111011101110;
20'b01010000110110101101: color_data = 12'b111011101110;
20'b01010000110110101110: color_data = 12'b111011101110;
20'b01010000110110101111: color_data = 12'b111011101110;
20'b01010000110110110000: color_data = 12'b111011101110;
20'b01010000110111001000: color_data = 12'b111011101110;
20'b01010000110111001001: color_data = 12'b111011101110;
20'b01010000110111001010: color_data = 12'b111011101110;
20'b01010000110111001011: color_data = 12'b111011101110;
20'b01010000110111001100: color_data = 12'b111011101110;
20'b01010000110111001101: color_data = 12'b111011101110;
20'b01010000110111001110: color_data = 12'b111011101110;
20'b01010000110111001111: color_data = 12'b111011101110;
20'b01010000110111010000: color_data = 12'b111011101110;
20'b01010000110111010001: color_data = 12'b111011101110;
20'b01010000110111010011: color_data = 12'b111011101110;
20'b01010000110111010100: color_data = 12'b111011101110;
20'b01010000110111010101: color_data = 12'b111011101110;
20'b01010000110111010110: color_data = 12'b111011101110;
20'b01010000110111010111: color_data = 12'b111011101110;
20'b01010000110111011000: color_data = 12'b111011101110;
20'b01010000110111011001: color_data = 12'b111011101110;
20'b01010000110111011010: color_data = 12'b111011101110;
20'b01010000110111011011: color_data = 12'b111011101110;
20'b01010000110111011100: color_data = 12'b111011101110;
20'b01010001000010100001: color_data = 12'b111011101110;
20'b01010001000010100010: color_data = 12'b111011101110;
20'b01010001000010100011: color_data = 12'b111011101110;
20'b01010001000010100100: color_data = 12'b111011101110;
20'b01010001000010100101: color_data = 12'b111011101110;
20'b01010001000010100110: color_data = 12'b111011101110;
20'b01010001000010100111: color_data = 12'b111011101110;
20'b01010001000010101000: color_data = 12'b111011101110;
20'b01010001000010101001: color_data = 12'b111011101110;
20'b01010001000010101010: color_data = 12'b111011101110;
20'b01010001000010101100: color_data = 12'b111011101110;
20'b01010001000010101101: color_data = 12'b111011101110;
20'b01010001000010101110: color_data = 12'b111011101110;
20'b01010001000010101111: color_data = 12'b111011101110;
20'b01010001000010110000: color_data = 12'b111011101110;
20'b01010001000010110001: color_data = 12'b111011101110;
20'b01010001000010110010: color_data = 12'b111011101110;
20'b01010001000010110011: color_data = 12'b111011101110;
20'b01010001000010110100: color_data = 12'b111011101110;
20'b01010001000010110101: color_data = 12'b111011101110;
20'b01010001000010110111: color_data = 12'b111011101110;
20'b01010001000010111000: color_data = 12'b111011101110;
20'b01010001000010111001: color_data = 12'b111011101110;
20'b01010001000010111010: color_data = 12'b111011101110;
20'b01010001000010111011: color_data = 12'b111011101110;
20'b01010001000010111100: color_data = 12'b111011101110;
20'b01010001000010111101: color_data = 12'b111011101110;
20'b01010001000010111110: color_data = 12'b111011101110;
20'b01010001000010111111: color_data = 12'b111011101110;
20'b01010001000011000000: color_data = 12'b111011101110;
20'b01010001000011000010: color_data = 12'b111011101110;
20'b01010001000011000011: color_data = 12'b111011101110;
20'b01010001000011000100: color_data = 12'b111011101110;
20'b01010001000011000101: color_data = 12'b111011101110;
20'b01010001000011000110: color_data = 12'b111011101110;
20'b01010001000011000111: color_data = 12'b111011101110;
20'b01010001000011001000: color_data = 12'b111011101110;
20'b01010001000011001001: color_data = 12'b111011101110;
20'b01010001000011001010: color_data = 12'b111011101110;
20'b01010001000011001011: color_data = 12'b111011101110;
20'b01010001000011001101: color_data = 12'b111011101110;
20'b01010001000011001110: color_data = 12'b111011101110;
20'b01010001000011001111: color_data = 12'b111011101110;
20'b01010001000011010000: color_data = 12'b111011101110;
20'b01010001000011010001: color_data = 12'b111011101110;
20'b01010001000011010010: color_data = 12'b111011101110;
20'b01010001000011010011: color_data = 12'b111011101110;
20'b01010001000011010100: color_data = 12'b111011101110;
20'b01010001000011010101: color_data = 12'b111011101110;
20'b01010001000011010110: color_data = 12'b111011101110;
20'b01010001000011111000: color_data = 12'b111011101110;
20'b01010001000011111001: color_data = 12'b111011101110;
20'b01010001000011111010: color_data = 12'b111011101110;
20'b01010001000011111011: color_data = 12'b111011101110;
20'b01010001000011111100: color_data = 12'b111011101110;
20'b01010001000011111101: color_data = 12'b111011101110;
20'b01010001000011111110: color_data = 12'b111011101110;
20'b01010001000011111111: color_data = 12'b111011101110;
20'b01010001000100000000: color_data = 12'b111011101110;
20'b01010001000100000001: color_data = 12'b111011101110;
20'b01010001000100000011: color_data = 12'b111011101110;
20'b01010001000100000100: color_data = 12'b111011101110;
20'b01010001000100000101: color_data = 12'b111011101110;
20'b01010001000100000110: color_data = 12'b111011101110;
20'b01010001000100000111: color_data = 12'b111011101110;
20'b01010001000100001000: color_data = 12'b111011101110;
20'b01010001000100001001: color_data = 12'b111011101110;
20'b01010001000100001010: color_data = 12'b111011101110;
20'b01010001000100001011: color_data = 12'b111011101110;
20'b01010001000100001100: color_data = 12'b111011101110;
20'b01010001000100001110: color_data = 12'b111011101110;
20'b01010001000100001111: color_data = 12'b111011101110;
20'b01010001000100010000: color_data = 12'b111011101110;
20'b01010001000100010001: color_data = 12'b111011101110;
20'b01010001000100010010: color_data = 12'b111011101110;
20'b01010001000100010011: color_data = 12'b111011101110;
20'b01010001000100010100: color_data = 12'b111011101110;
20'b01010001000100010101: color_data = 12'b111011101110;
20'b01010001000100010110: color_data = 12'b111011101110;
20'b01010001000100010111: color_data = 12'b111011101110;
20'b01010001000100011001: color_data = 12'b111011101110;
20'b01010001000100011010: color_data = 12'b111011101110;
20'b01010001000100011011: color_data = 12'b111011101110;
20'b01010001000100011100: color_data = 12'b111011101110;
20'b01010001000100011101: color_data = 12'b111011101110;
20'b01010001000100011110: color_data = 12'b111011101110;
20'b01010001000100011111: color_data = 12'b111011101110;
20'b01010001000100100000: color_data = 12'b111011101110;
20'b01010001000100100001: color_data = 12'b111011101110;
20'b01010001000100100010: color_data = 12'b111011101110;
20'b01010001000100100100: color_data = 12'b111011101110;
20'b01010001000100100101: color_data = 12'b111011101110;
20'b01010001000100100110: color_data = 12'b111011101110;
20'b01010001000100100111: color_data = 12'b111011101110;
20'b01010001000100101000: color_data = 12'b111011101110;
20'b01010001000100101001: color_data = 12'b111011101110;
20'b01010001000100101010: color_data = 12'b111011101110;
20'b01010001000100101011: color_data = 12'b111011101110;
20'b01010001000100101100: color_data = 12'b111011101110;
20'b01010001000100101101: color_data = 12'b111011101110;
20'b01010001000101000100: color_data = 12'b111011101110;
20'b01010001000101000101: color_data = 12'b111011101110;
20'b01010001000101000110: color_data = 12'b111011101110;
20'b01010001000101000111: color_data = 12'b111011101110;
20'b01010001000101001000: color_data = 12'b111011101110;
20'b01010001000101001001: color_data = 12'b111011101110;
20'b01010001000101001010: color_data = 12'b111011101110;
20'b01010001000101001011: color_data = 12'b111011101110;
20'b01010001000101001100: color_data = 12'b111011101110;
20'b01010001000101001101: color_data = 12'b111011101110;
20'b01010001000101001111: color_data = 12'b111011101110;
20'b01010001000101010000: color_data = 12'b111011101110;
20'b01010001000101010001: color_data = 12'b111011101110;
20'b01010001000101010010: color_data = 12'b111011101110;
20'b01010001000101010011: color_data = 12'b111011101110;
20'b01010001000101010100: color_data = 12'b111011101110;
20'b01010001000101010101: color_data = 12'b111011101110;
20'b01010001000101010110: color_data = 12'b111011101110;
20'b01010001000101010111: color_data = 12'b111011101110;
20'b01010001000101011000: color_data = 12'b111011101110;
20'b01010001000101011010: color_data = 12'b111011101110;
20'b01010001000101011011: color_data = 12'b111011101110;
20'b01010001000101011100: color_data = 12'b111011101110;
20'b01010001000101011101: color_data = 12'b111011101110;
20'b01010001000101011110: color_data = 12'b111011101110;
20'b01010001000101011111: color_data = 12'b111011101110;
20'b01010001000101100000: color_data = 12'b111011101110;
20'b01010001000101100001: color_data = 12'b111011101110;
20'b01010001000101100010: color_data = 12'b111011101110;
20'b01010001000101100011: color_data = 12'b111011101110;
20'b01010001000101100101: color_data = 12'b111011101110;
20'b01010001000101100110: color_data = 12'b111011101110;
20'b01010001000101100111: color_data = 12'b111011101110;
20'b01010001000101101000: color_data = 12'b111011101110;
20'b01010001000101101001: color_data = 12'b111011101110;
20'b01010001000101101010: color_data = 12'b111011101110;
20'b01010001000101101011: color_data = 12'b111011101110;
20'b01010001000101101100: color_data = 12'b111011101110;
20'b01010001000101101101: color_data = 12'b111011101110;
20'b01010001000101101110: color_data = 12'b111011101110;
20'b01010001000101110000: color_data = 12'b111011101110;
20'b01010001000101110001: color_data = 12'b111011101110;
20'b01010001000101110010: color_data = 12'b111011101110;
20'b01010001000101110011: color_data = 12'b111011101110;
20'b01010001000101110100: color_data = 12'b111011101110;
20'b01010001000101110101: color_data = 12'b111011101110;
20'b01010001000101110110: color_data = 12'b111011101110;
20'b01010001000101110111: color_data = 12'b111011101110;
20'b01010001000101111000: color_data = 12'b111011101110;
20'b01010001000101111001: color_data = 12'b111011101110;
20'b01010001000101111011: color_data = 12'b111011101110;
20'b01010001000101111100: color_data = 12'b111011101110;
20'b01010001000101111101: color_data = 12'b111011101110;
20'b01010001000101111110: color_data = 12'b111011101110;
20'b01010001000101111111: color_data = 12'b111011101110;
20'b01010001000110000000: color_data = 12'b111011101110;
20'b01010001000110000001: color_data = 12'b111011101110;
20'b01010001000110000010: color_data = 12'b111011101110;
20'b01010001000110000011: color_data = 12'b111011101110;
20'b01010001000110000100: color_data = 12'b111011101110;
20'b01010001000110000110: color_data = 12'b111011101110;
20'b01010001000110000111: color_data = 12'b111011101110;
20'b01010001000110001000: color_data = 12'b111011101110;
20'b01010001000110001001: color_data = 12'b111011101110;
20'b01010001000110001010: color_data = 12'b111011101110;
20'b01010001000110001011: color_data = 12'b111011101110;
20'b01010001000110001100: color_data = 12'b111011101110;
20'b01010001000110001101: color_data = 12'b111011101110;
20'b01010001000110001110: color_data = 12'b111011101110;
20'b01010001000110001111: color_data = 12'b111011101110;
20'b01010001000110011100: color_data = 12'b111011101110;
20'b01010001000110011101: color_data = 12'b111011101110;
20'b01010001000110011110: color_data = 12'b111011101110;
20'b01010001000110011111: color_data = 12'b111011101110;
20'b01010001000110100000: color_data = 12'b111011101110;
20'b01010001000110100001: color_data = 12'b111011101110;
20'b01010001000110100010: color_data = 12'b111011101110;
20'b01010001000110100011: color_data = 12'b111011101110;
20'b01010001000110100100: color_data = 12'b111011101110;
20'b01010001000110100101: color_data = 12'b111011101110;
20'b01010001000110100111: color_data = 12'b111011101110;
20'b01010001000110101000: color_data = 12'b111011101110;
20'b01010001000110101001: color_data = 12'b111011101110;
20'b01010001000110101010: color_data = 12'b111011101110;
20'b01010001000110101011: color_data = 12'b111011101110;
20'b01010001000110101100: color_data = 12'b111011101110;
20'b01010001000110101101: color_data = 12'b111011101110;
20'b01010001000110101110: color_data = 12'b111011101110;
20'b01010001000110101111: color_data = 12'b111011101110;
20'b01010001000110110000: color_data = 12'b111011101110;
20'b01010001000111001000: color_data = 12'b111011101110;
20'b01010001000111001001: color_data = 12'b111011101110;
20'b01010001000111001010: color_data = 12'b111011101110;
20'b01010001000111001011: color_data = 12'b111011101110;
20'b01010001000111001100: color_data = 12'b111011101110;
20'b01010001000111001101: color_data = 12'b111011101110;
20'b01010001000111001110: color_data = 12'b111011101110;
20'b01010001000111001111: color_data = 12'b111011101110;
20'b01010001000111010000: color_data = 12'b111011101110;
20'b01010001000111010001: color_data = 12'b111011101110;
20'b01010001000111010011: color_data = 12'b111011101110;
20'b01010001000111010100: color_data = 12'b111011101110;
20'b01010001000111010101: color_data = 12'b111011101110;
20'b01010001000111010110: color_data = 12'b111011101110;
20'b01010001000111010111: color_data = 12'b111011101110;
20'b01010001000111011000: color_data = 12'b111011101110;
20'b01010001000111011001: color_data = 12'b111011101110;
20'b01010001000111011010: color_data = 12'b111011101110;
20'b01010001000111011011: color_data = 12'b111011101110;
20'b01010001000111011100: color_data = 12'b111011101110;
20'b01010001010010100001: color_data = 12'b111011101110;
20'b01010001010010100010: color_data = 12'b111011101110;
20'b01010001010010100011: color_data = 12'b111011101110;
20'b01010001010010100100: color_data = 12'b111011101110;
20'b01010001010010100101: color_data = 12'b111011101110;
20'b01010001010010100110: color_data = 12'b111011101110;
20'b01010001010010100111: color_data = 12'b111011101110;
20'b01010001010010101000: color_data = 12'b111011101110;
20'b01010001010010101001: color_data = 12'b111011101110;
20'b01010001010010101010: color_data = 12'b111011101110;
20'b01010001010010101100: color_data = 12'b111011101110;
20'b01010001010010101101: color_data = 12'b111011101110;
20'b01010001010010101110: color_data = 12'b111011101110;
20'b01010001010010101111: color_data = 12'b111011101110;
20'b01010001010010110000: color_data = 12'b111011101110;
20'b01010001010010110001: color_data = 12'b111011101110;
20'b01010001010010110010: color_data = 12'b111011101110;
20'b01010001010010110011: color_data = 12'b111011101110;
20'b01010001010010110100: color_data = 12'b111011101110;
20'b01010001010010110101: color_data = 12'b111011101110;
20'b01010001010010110111: color_data = 12'b111011101110;
20'b01010001010010111000: color_data = 12'b111011101110;
20'b01010001010010111001: color_data = 12'b111011101110;
20'b01010001010010111010: color_data = 12'b111011101110;
20'b01010001010010111011: color_data = 12'b111011101110;
20'b01010001010010111100: color_data = 12'b111011101110;
20'b01010001010010111101: color_data = 12'b111011101110;
20'b01010001010010111110: color_data = 12'b111011101110;
20'b01010001010010111111: color_data = 12'b111011101110;
20'b01010001010011000000: color_data = 12'b111011101110;
20'b01010001010011000010: color_data = 12'b111011101110;
20'b01010001010011000011: color_data = 12'b111011101110;
20'b01010001010011000100: color_data = 12'b111011101110;
20'b01010001010011000101: color_data = 12'b111011101110;
20'b01010001010011000110: color_data = 12'b111011101110;
20'b01010001010011000111: color_data = 12'b111011101110;
20'b01010001010011001000: color_data = 12'b111011101110;
20'b01010001010011001001: color_data = 12'b111011101110;
20'b01010001010011001010: color_data = 12'b111011101110;
20'b01010001010011001011: color_data = 12'b111011101110;
20'b01010001010011001101: color_data = 12'b111011101110;
20'b01010001010011001110: color_data = 12'b111011101110;
20'b01010001010011001111: color_data = 12'b111011101110;
20'b01010001010011010000: color_data = 12'b111011101110;
20'b01010001010011010001: color_data = 12'b111011101110;
20'b01010001010011010010: color_data = 12'b111011101110;
20'b01010001010011010011: color_data = 12'b111011101110;
20'b01010001010011010100: color_data = 12'b111011101110;
20'b01010001010011010101: color_data = 12'b111011101110;
20'b01010001010011010110: color_data = 12'b111011101110;
20'b01010001010011111000: color_data = 12'b111011101110;
20'b01010001010011111001: color_data = 12'b111011101110;
20'b01010001010011111010: color_data = 12'b111011101110;
20'b01010001010011111011: color_data = 12'b111011101110;
20'b01010001010011111100: color_data = 12'b111011101110;
20'b01010001010011111101: color_data = 12'b111011101110;
20'b01010001010011111110: color_data = 12'b111011101110;
20'b01010001010011111111: color_data = 12'b111011101110;
20'b01010001010100000000: color_data = 12'b111011101110;
20'b01010001010100000001: color_data = 12'b111011101110;
20'b01010001010100000011: color_data = 12'b111011101110;
20'b01010001010100000100: color_data = 12'b111011101110;
20'b01010001010100000101: color_data = 12'b111011101110;
20'b01010001010100000110: color_data = 12'b111011101110;
20'b01010001010100000111: color_data = 12'b111011101110;
20'b01010001010100001000: color_data = 12'b111011101110;
20'b01010001010100001001: color_data = 12'b111011101110;
20'b01010001010100001010: color_data = 12'b111011101110;
20'b01010001010100001011: color_data = 12'b111011101110;
20'b01010001010100001100: color_data = 12'b111011101110;
20'b01010001010100001110: color_data = 12'b111011101110;
20'b01010001010100001111: color_data = 12'b111011101110;
20'b01010001010100010000: color_data = 12'b111011101110;
20'b01010001010100010001: color_data = 12'b111011101110;
20'b01010001010100010010: color_data = 12'b111011101110;
20'b01010001010100010011: color_data = 12'b111011101110;
20'b01010001010100010100: color_data = 12'b111011101110;
20'b01010001010100010101: color_data = 12'b111011101110;
20'b01010001010100010110: color_data = 12'b111011101110;
20'b01010001010100010111: color_data = 12'b111011101110;
20'b01010001010100011001: color_data = 12'b111011101110;
20'b01010001010100011010: color_data = 12'b111011101110;
20'b01010001010100011011: color_data = 12'b111011101110;
20'b01010001010100011100: color_data = 12'b111011101110;
20'b01010001010100011101: color_data = 12'b111011101110;
20'b01010001010100011110: color_data = 12'b111011101110;
20'b01010001010100011111: color_data = 12'b111011101110;
20'b01010001010100100000: color_data = 12'b111011101110;
20'b01010001010100100001: color_data = 12'b111011101110;
20'b01010001010100100010: color_data = 12'b111011101110;
20'b01010001010100100100: color_data = 12'b111011101110;
20'b01010001010100100101: color_data = 12'b111011101110;
20'b01010001010100100110: color_data = 12'b111011101110;
20'b01010001010100100111: color_data = 12'b111011101110;
20'b01010001010100101000: color_data = 12'b111011101110;
20'b01010001010100101001: color_data = 12'b111011101110;
20'b01010001010100101010: color_data = 12'b111011101110;
20'b01010001010100101011: color_data = 12'b111011101110;
20'b01010001010100101100: color_data = 12'b111011101110;
20'b01010001010100101101: color_data = 12'b111011101110;
20'b01010001010101000100: color_data = 12'b111011101110;
20'b01010001010101000101: color_data = 12'b111011101110;
20'b01010001010101000110: color_data = 12'b111011101110;
20'b01010001010101000111: color_data = 12'b111011101110;
20'b01010001010101001000: color_data = 12'b111011101110;
20'b01010001010101001001: color_data = 12'b111011101110;
20'b01010001010101001010: color_data = 12'b111011101110;
20'b01010001010101001011: color_data = 12'b111011101110;
20'b01010001010101001100: color_data = 12'b111011101110;
20'b01010001010101001101: color_data = 12'b111011101110;
20'b01010001010101001111: color_data = 12'b111011101110;
20'b01010001010101010000: color_data = 12'b111011101110;
20'b01010001010101010001: color_data = 12'b111011101110;
20'b01010001010101010010: color_data = 12'b111011101110;
20'b01010001010101010011: color_data = 12'b111011101110;
20'b01010001010101010100: color_data = 12'b111011101110;
20'b01010001010101010101: color_data = 12'b111011101110;
20'b01010001010101010110: color_data = 12'b111011101110;
20'b01010001010101010111: color_data = 12'b111011101110;
20'b01010001010101011000: color_data = 12'b111011101110;
20'b01010001010101011010: color_data = 12'b111011101110;
20'b01010001010101011011: color_data = 12'b111011101110;
20'b01010001010101011100: color_data = 12'b111011101110;
20'b01010001010101011101: color_data = 12'b111011101110;
20'b01010001010101011110: color_data = 12'b111011101110;
20'b01010001010101011111: color_data = 12'b111011101110;
20'b01010001010101100000: color_data = 12'b111011101110;
20'b01010001010101100001: color_data = 12'b111011101110;
20'b01010001010101100010: color_data = 12'b111011101110;
20'b01010001010101100011: color_data = 12'b111011101110;
20'b01010001010101100101: color_data = 12'b111011101110;
20'b01010001010101100110: color_data = 12'b111011101110;
20'b01010001010101100111: color_data = 12'b111011101110;
20'b01010001010101101000: color_data = 12'b111011101110;
20'b01010001010101101001: color_data = 12'b111011101110;
20'b01010001010101101010: color_data = 12'b111011101110;
20'b01010001010101101011: color_data = 12'b111011101110;
20'b01010001010101101100: color_data = 12'b111011101110;
20'b01010001010101101101: color_data = 12'b111011101110;
20'b01010001010101101110: color_data = 12'b111011101110;
20'b01010001010101110000: color_data = 12'b111011101110;
20'b01010001010101110001: color_data = 12'b111011101110;
20'b01010001010101110010: color_data = 12'b111011101110;
20'b01010001010101110011: color_data = 12'b111011101110;
20'b01010001010101110100: color_data = 12'b111011101110;
20'b01010001010101110101: color_data = 12'b111011101110;
20'b01010001010101110110: color_data = 12'b111011101110;
20'b01010001010101110111: color_data = 12'b111011101110;
20'b01010001010101111000: color_data = 12'b111011101110;
20'b01010001010101111001: color_data = 12'b111011101110;
20'b01010001010101111011: color_data = 12'b111011101110;
20'b01010001010101111100: color_data = 12'b111011101110;
20'b01010001010101111101: color_data = 12'b111011101110;
20'b01010001010101111110: color_data = 12'b111011101110;
20'b01010001010101111111: color_data = 12'b111011101110;
20'b01010001010110000000: color_data = 12'b111011101110;
20'b01010001010110000001: color_data = 12'b111011101110;
20'b01010001010110000010: color_data = 12'b111011101110;
20'b01010001010110000011: color_data = 12'b111011101110;
20'b01010001010110000100: color_data = 12'b111011101110;
20'b01010001010110000110: color_data = 12'b111011101110;
20'b01010001010110000111: color_data = 12'b111011101110;
20'b01010001010110001000: color_data = 12'b111011101110;
20'b01010001010110001001: color_data = 12'b111011101110;
20'b01010001010110001010: color_data = 12'b111011101110;
20'b01010001010110001011: color_data = 12'b111011101110;
20'b01010001010110001100: color_data = 12'b111011101110;
20'b01010001010110001101: color_data = 12'b111011101110;
20'b01010001010110001110: color_data = 12'b111011101110;
20'b01010001010110001111: color_data = 12'b111011101110;
20'b01010001010110011100: color_data = 12'b111011101110;
20'b01010001010110011101: color_data = 12'b111011101110;
20'b01010001010110011110: color_data = 12'b111011101110;
20'b01010001010110011111: color_data = 12'b111011101110;
20'b01010001010110100000: color_data = 12'b111011101110;
20'b01010001010110100001: color_data = 12'b111011101110;
20'b01010001010110100010: color_data = 12'b111011101110;
20'b01010001010110100011: color_data = 12'b111011101110;
20'b01010001010110100100: color_data = 12'b111011101110;
20'b01010001010110100101: color_data = 12'b111011101110;
20'b01010001010110100111: color_data = 12'b111011101110;
20'b01010001010110101000: color_data = 12'b111011101110;
20'b01010001010110101001: color_data = 12'b111011101110;
20'b01010001010110101010: color_data = 12'b111011101110;
20'b01010001010110101011: color_data = 12'b111011101110;
20'b01010001010110101100: color_data = 12'b111011101110;
20'b01010001010110101101: color_data = 12'b111011101110;
20'b01010001010110101110: color_data = 12'b111011101110;
20'b01010001010110101111: color_data = 12'b111011101110;
20'b01010001010110110000: color_data = 12'b111011101110;
20'b01010001010111001000: color_data = 12'b111011101110;
20'b01010001010111001001: color_data = 12'b111011101110;
20'b01010001010111001010: color_data = 12'b111011101110;
20'b01010001010111001011: color_data = 12'b111011101110;
20'b01010001010111001100: color_data = 12'b111011101110;
20'b01010001010111001101: color_data = 12'b111011101110;
20'b01010001010111001110: color_data = 12'b111011101110;
20'b01010001010111001111: color_data = 12'b111011101110;
20'b01010001010111010000: color_data = 12'b111011101110;
20'b01010001010111010001: color_data = 12'b111011101110;
20'b01010001010111010011: color_data = 12'b111011101110;
20'b01010001010111010100: color_data = 12'b111011101110;
20'b01010001010111010101: color_data = 12'b111011101110;
20'b01010001010111010110: color_data = 12'b111011101110;
20'b01010001010111010111: color_data = 12'b111011101110;
20'b01010001010111011000: color_data = 12'b111011101110;
20'b01010001010111011001: color_data = 12'b111011101110;
20'b01010001010111011010: color_data = 12'b111011101110;
20'b01010001010111011011: color_data = 12'b111011101110;
20'b01010001010111011100: color_data = 12'b111011101110;
20'b01010001100010100001: color_data = 12'b111011101110;
20'b01010001100010100010: color_data = 12'b111011101110;
20'b01010001100010100011: color_data = 12'b111011101110;
20'b01010001100010100100: color_data = 12'b111011101110;
20'b01010001100010100101: color_data = 12'b111011101110;
20'b01010001100010100110: color_data = 12'b111011101110;
20'b01010001100010100111: color_data = 12'b111011101110;
20'b01010001100010101000: color_data = 12'b111011101110;
20'b01010001100010101001: color_data = 12'b111011101110;
20'b01010001100010101010: color_data = 12'b111011101110;
20'b01010001100010101100: color_data = 12'b111011101110;
20'b01010001100010101101: color_data = 12'b111011101110;
20'b01010001100010101110: color_data = 12'b111011101110;
20'b01010001100010101111: color_data = 12'b111011101110;
20'b01010001100010110000: color_data = 12'b111011101110;
20'b01010001100010110001: color_data = 12'b111011101110;
20'b01010001100010110010: color_data = 12'b111011101110;
20'b01010001100010110011: color_data = 12'b111011101110;
20'b01010001100010110100: color_data = 12'b111011101110;
20'b01010001100010110101: color_data = 12'b111011101110;
20'b01010001100010110111: color_data = 12'b111011101110;
20'b01010001100010111000: color_data = 12'b111011101110;
20'b01010001100010111001: color_data = 12'b111011101110;
20'b01010001100010111010: color_data = 12'b111011101110;
20'b01010001100010111011: color_data = 12'b111011101110;
20'b01010001100010111100: color_data = 12'b111011101110;
20'b01010001100010111101: color_data = 12'b111011101110;
20'b01010001100010111110: color_data = 12'b111011101110;
20'b01010001100010111111: color_data = 12'b111011101110;
20'b01010001100011000000: color_data = 12'b111011101110;
20'b01010001100011000010: color_data = 12'b111011101110;
20'b01010001100011000011: color_data = 12'b111011101110;
20'b01010001100011000100: color_data = 12'b111011101110;
20'b01010001100011000101: color_data = 12'b111011101110;
20'b01010001100011000110: color_data = 12'b111011101110;
20'b01010001100011000111: color_data = 12'b111011101110;
20'b01010001100011001000: color_data = 12'b111011101110;
20'b01010001100011001001: color_data = 12'b111011101110;
20'b01010001100011001010: color_data = 12'b111011101110;
20'b01010001100011001011: color_data = 12'b111011101110;
20'b01010001100011001101: color_data = 12'b111011101110;
20'b01010001100011001110: color_data = 12'b111011101110;
20'b01010001100011001111: color_data = 12'b111011101110;
20'b01010001100011010000: color_data = 12'b111011101110;
20'b01010001100011010001: color_data = 12'b111011101110;
20'b01010001100011010010: color_data = 12'b111011101110;
20'b01010001100011010011: color_data = 12'b111011101110;
20'b01010001100011010100: color_data = 12'b111011101110;
20'b01010001100011010101: color_data = 12'b111011101110;
20'b01010001100011010110: color_data = 12'b111011101110;
20'b01010001100011111000: color_data = 12'b111011101110;
20'b01010001100011111001: color_data = 12'b111011101110;
20'b01010001100011111010: color_data = 12'b111011101110;
20'b01010001100011111011: color_data = 12'b111011101110;
20'b01010001100011111100: color_data = 12'b111011101110;
20'b01010001100011111101: color_data = 12'b111011101110;
20'b01010001100011111110: color_data = 12'b111011101110;
20'b01010001100011111111: color_data = 12'b111011101110;
20'b01010001100100000000: color_data = 12'b111011101110;
20'b01010001100100000001: color_data = 12'b111011101110;
20'b01010001100100000011: color_data = 12'b111011101110;
20'b01010001100100000100: color_data = 12'b111011101110;
20'b01010001100100000101: color_data = 12'b111011101110;
20'b01010001100100000110: color_data = 12'b111011101110;
20'b01010001100100000111: color_data = 12'b111011101110;
20'b01010001100100001000: color_data = 12'b111011101110;
20'b01010001100100001001: color_data = 12'b111011101110;
20'b01010001100100001010: color_data = 12'b111011101110;
20'b01010001100100001011: color_data = 12'b111011101110;
20'b01010001100100001100: color_data = 12'b111011101110;
20'b01010001100100001110: color_data = 12'b111011101110;
20'b01010001100100001111: color_data = 12'b111011101110;
20'b01010001100100010000: color_data = 12'b111011101110;
20'b01010001100100010001: color_data = 12'b111011101110;
20'b01010001100100010010: color_data = 12'b111011101110;
20'b01010001100100010011: color_data = 12'b111011101110;
20'b01010001100100010100: color_data = 12'b111011101110;
20'b01010001100100010101: color_data = 12'b111011101110;
20'b01010001100100010110: color_data = 12'b111011101110;
20'b01010001100100010111: color_data = 12'b111011101110;
20'b01010001100100011001: color_data = 12'b111011101110;
20'b01010001100100011010: color_data = 12'b111011101110;
20'b01010001100100011011: color_data = 12'b111011101110;
20'b01010001100100011100: color_data = 12'b111011101110;
20'b01010001100100011101: color_data = 12'b111011101110;
20'b01010001100100011110: color_data = 12'b111011101110;
20'b01010001100100011111: color_data = 12'b111011101110;
20'b01010001100100100000: color_data = 12'b111011101110;
20'b01010001100100100001: color_data = 12'b111011101110;
20'b01010001100100100010: color_data = 12'b111011101110;
20'b01010001100100100100: color_data = 12'b111011101110;
20'b01010001100100100101: color_data = 12'b111011101110;
20'b01010001100100100110: color_data = 12'b111011101110;
20'b01010001100100100111: color_data = 12'b111011101110;
20'b01010001100100101000: color_data = 12'b111011101110;
20'b01010001100100101001: color_data = 12'b111011101110;
20'b01010001100100101010: color_data = 12'b111011101110;
20'b01010001100100101011: color_data = 12'b111011101110;
20'b01010001100100101100: color_data = 12'b111011101110;
20'b01010001100100101101: color_data = 12'b111011101110;
20'b01010001100101000100: color_data = 12'b111011101110;
20'b01010001100101000101: color_data = 12'b111011101110;
20'b01010001100101000110: color_data = 12'b111011101110;
20'b01010001100101000111: color_data = 12'b111011101110;
20'b01010001100101001000: color_data = 12'b111011101110;
20'b01010001100101001001: color_data = 12'b111011101110;
20'b01010001100101001010: color_data = 12'b111011101110;
20'b01010001100101001011: color_data = 12'b111011101110;
20'b01010001100101001100: color_data = 12'b111011101110;
20'b01010001100101001101: color_data = 12'b111011101110;
20'b01010001100101001111: color_data = 12'b111011101110;
20'b01010001100101010000: color_data = 12'b111011101110;
20'b01010001100101010001: color_data = 12'b111011101110;
20'b01010001100101010010: color_data = 12'b111011101110;
20'b01010001100101010011: color_data = 12'b111011101110;
20'b01010001100101010100: color_data = 12'b111011101110;
20'b01010001100101010101: color_data = 12'b111011101110;
20'b01010001100101010110: color_data = 12'b111011101110;
20'b01010001100101010111: color_data = 12'b111011101110;
20'b01010001100101011000: color_data = 12'b111011101110;
20'b01010001100101011010: color_data = 12'b111011101110;
20'b01010001100101011011: color_data = 12'b111011101110;
20'b01010001100101011100: color_data = 12'b111011101110;
20'b01010001100101011101: color_data = 12'b111011101110;
20'b01010001100101011110: color_data = 12'b111011101110;
20'b01010001100101011111: color_data = 12'b111011101110;
20'b01010001100101100000: color_data = 12'b111011101110;
20'b01010001100101100001: color_data = 12'b111011101110;
20'b01010001100101100010: color_data = 12'b111011101110;
20'b01010001100101100011: color_data = 12'b111011101110;
20'b01010001100101100101: color_data = 12'b111011101110;
20'b01010001100101100110: color_data = 12'b111011101110;
20'b01010001100101100111: color_data = 12'b111011101110;
20'b01010001100101101000: color_data = 12'b111011101110;
20'b01010001100101101001: color_data = 12'b111011101110;
20'b01010001100101101010: color_data = 12'b111011101110;
20'b01010001100101101011: color_data = 12'b111011101110;
20'b01010001100101101100: color_data = 12'b111011101110;
20'b01010001100101101101: color_data = 12'b111011101110;
20'b01010001100101101110: color_data = 12'b111011101110;
20'b01010001100101110000: color_data = 12'b111011101110;
20'b01010001100101110001: color_data = 12'b111011101110;
20'b01010001100101110010: color_data = 12'b111011101110;
20'b01010001100101110011: color_data = 12'b111011101110;
20'b01010001100101110100: color_data = 12'b111011101110;
20'b01010001100101110101: color_data = 12'b111011101110;
20'b01010001100101110110: color_data = 12'b111011101110;
20'b01010001100101110111: color_data = 12'b111011101110;
20'b01010001100101111000: color_data = 12'b111011101110;
20'b01010001100101111001: color_data = 12'b111011101110;
20'b01010001100101111011: color_data = 12'b111011101110;
20'b01010001100101111100: color_data = 12'b111011101110;
20'b01010001100101111101: color_data = 12'b111011101110;
20'b01010001100101111110: color_data = 12'b111011101110;
20'b01010001100101111111: color_data = 12'b111011101110;
20'b01010001100110000000: color_data = 12'b111011101110;
20'b01010001100110000001: color_data = 12'b111011101110;
20'b01010001100110000010: color_data = 12'b111011101110;
20'b01010001100110000011: color_data = 12'b111011101110;
20'b01010001100110000100: color_data = 12'b111011101110;
20'b01010001100110000110: color_data = 12'b111011101110;
20'b01010001100110000111: color_data = 12'b111011101110;
20'b01010001100110001000: color_data = 12'b111011101110;
20'b01010001100110001001: color_data = 12'b111011101110;
20'b01010001100110001010: color_data = 12'b111011101110;
20'b01010001100110001011: color_data = 12'b111011101110;
20'b01010001100110001100: color_data = 12'b111011101110;
20'b01010001100110001101: color_data = 12'b111011101110;
20'b01010001100110001110: color_data = 12'b111011101110;
20'b01010001100110001111: color_data = 12'b111011101110;
20'b01010001100110011100: color_data = 12'b111011101110;
20'b01010001100110011101: color_data = 12'b111011101110;
20'b01010001100110011110: color_data = 12'b111011101110;
20'b01010001100110011111: color_data = 12'b111011101110;
20'b01010001100110100000: color_data = 12'b111011101110;
20'b01010001100110100001: color_data = 12'b111011101110;
20'b01010001100110100010: color_data = 12'b111011101110;
20'b01010001100110100011: color_data = 12'b111011101110;
20'b01010001100110100100: color_data = 12'b111011101110;
20'b01010001100110100101: color_data = 12'b111011101110;
20'b01010001100110100111: color_data = 12'b111011101110;
20'b01010001100110101000: color_data = 12'b111011101110;
20'b01010001100110101001: color_data = 12'b111011101110;
20'b01010001100110101010: color_data = 12'b111011101110;
20'b01010001100110101011: color_data = 12'b111011101110;
20'b01010001100110101100: color_data = 12'b111011101110;
20'b01010001100110101101: color_data = 12'b111011101110;
20'b01010001100110101110: color_data = 12'b111011101110;
20'b01010001100110101111: color_data = 12'b111011101110;
20'b01010001100110110000: color_data = 12'b111011101110;
20'b01010001100111001000: color_data = 12'b111011101110;
20'b01010001100111001001: color_data = 12'b111011101110;
20'b01010001100111001010: color_data = 12'b111011101110;
20'b01010001100111001011: color_data = 12'b111011101110;
20'b01010001100111001100: color_data = 12'b111011101110;
20'b01010001100111001101: color_data = 12'b111011101110;
20'b01010001100111001110: color_data = 12'b111011101110;
20'b01010001100111001111: color_data = 12'b111011101110;
20'b01010001100111010000: color_data = 12'b111011101110;
20'b01010001100111010001: color_data = 12'b111011101110;
20'b01010001100111010011: color_data = 12'b111011101110;
20'b01010001100111010100: color_data = 12'b111011101110;
20'b01010001100111010101: color_data = 12'b111011101110;
20'b01010001100111010110: color_data = 12'b111011101110;
20'b01010001100111010111: color_data = 12'b111011101110;
20'b01010001100111011000: color_data = 12'b111011101110;
20'b01010001100111011001: color_data = 12'b111011101110;
20'b01010001100111011010: color_data = 12'b111011101110;
20'b01010001100111011011: color_data = 12'b111011101110;
20'b01010001100111011100: color_data = 12'b111011101110;
20'b01010001110010100001: color_data = 12'b111011101110;
20'b01010001110010100010: color_data = 12'b111011101110;
20'b01010001110010100011: color_data = 12'b111011101110;
20'b01010001110010100100: color_data = 12'b111011101110;
20'b01010001110010100101: color_data = 12'b111011101110;
20'b01010001110010100110: color_data = 12'b111011101110;
20'b01010001110010100111: color_data = 12'b111011101110;
20'b01010001110010101000: color_data = 12'b111011101110;
20'b01010001110010101001: color_data = 12'b111011101110;
20'b01010001110010101010: color_data = 12'b111011101110;
20'b01010001110010101100: color_data = 12'b111011101110;
20'b01010001110010101101: color_data = 12'b111011101110;
20'b01010001110010101110: color_data = 12'b111011101110;
20'b01010001110010101111: color_data = 12'b111011101110;
20'b01010001110010110000: color_data = 12'b111011101110;
20'b01010001110010110001: color_data = 12'b111011101110;
20'b01010001110010110010: color_data = 12'b111011101110;
20'b01010001110010110011: color_data = 12'b111011101110;
20'b01010001110010110100: color_data = 12'b111011101110;
20'b01010001110010110101: color_data = 12'b111011101110;
20'b01010001110010110111: color_data = 12'b111011101110;
20'b01010001110010111000: color_data = 12'b111011101110;
20'b01010001110010111001: color_data = 12'b111011101110;
20'b01010001110010111010: color_data = 12'b111011101110;
20'b01010001110010111011: color_data = 12'b111011101110;
20'b01010001110010111100: color_data = 12'b111011101110;
20'b01010001110010111101: color_data = 12'b111011101110;
20'b01010001110010111110: color_data = 12'b111011101110;
20'b01010001110010111111: color_data = 12'b111011101110;
20'b01010001110011000000: color_data = 12'b111011101110;
20'b01010001110011000010: color_data = 12'b111011101110;
20'b01010001110011000011: color_data = 12'b111011101110;
20'b01010001110011000100: color_data = 12'b111011101110;
20'b01010001110011000101: color_data = 12'b111011101110;
20'b01010001110011000110: color_data = 12'b111011101110;
20'b01010001110011000111: color_data = 12'b111011101110;
20'b01010001110011001000: color_data = 12'b111011101110;
20'b01010001110011001001: color_data = 12'b111011101110;
20'b01010001110011001010: color_data = 12'b111011101110;
20'b01010001110011001011: color_data = 12'b111011101110;
20'b01010001110011001101: color_data = 12'b111011101110;
20'b01010001110011001110: color_data = 12'b111011101110;
20'b01010001110011001111: color_data = 12'b111011101110;
20'b01010001110011010000: color_data = 12'b111011101110;
20'b01010001110011010001: color_data = 12'b111011101110;
20'b01010001110011010010: color_data = 12'b111011101110;
20'b01010001110011010011: color_data = 12'b111011101110;
20'b01010001110011010100: color_data = 12'b111011101110;
20'b01010001110011010101: color_data = 12'b111011101110;
20'b01010001110011010110: color_data = 12'b111011101110;
20'b01010001110011111000: color_data = 12'b111011101110;
20'b01010001110011111001: color_data = 12'b111011101110;
20'b01010001110011111010: color_data = 12'b111011101110;
20'b01010001110011111011: color_data = 12'b111011101110;
20'b01010001110011111100: color_data = 12'b111011101110;
20'b01010001110011111101: color_data = 12'b111011101110;
20'b01010001110011111110: color_data = 12'b111011101110;
20'b01010001110011111111: color_data = 12'b111011101110;
20'b01010001110100000000: color_data = 12'b111011101110;
20'b01010001110100000001: color_data = 12'b111011101110;
20'b01010001110100000011: color_data = 12'b111011101110;
20'b01010001110100000100: color_data = 12'b111011101110;
20'b01010001110100000101: color_data = 12'b111011101110;
20'b01010001110100000110: color_data = 12'b111011101110;
20'b01010001110100000111: color_data = 12'b111011101110;
20'b01010001110100001000: color_data = 12'b111011101110;
20'b01010001110100001001: color_data = 12'b111011101110;
20'b01010001110100001010: color_data = 12'b111011101110;
20'b01010001110100001011: color_data = 12'b111011101110;
20'b01010001110100001100: color_data = 12'b111011101110;
20'b01010001110100001110: color_data = 12'b111011101110;
20'b01010001110100001111: color_data = 12'b111011101110;
20'b01010001110100010000: color_data = 12'b111011101110;
20'b01010001110100010001: color_data = 12'b111011101110;
20'b01010001110100010010: color_data = 12'b111011101110;
20'b01010001110100010011: color_data = 12'b111011101110;
20'b01010001110100010100: color_data = 12'b111011101110;
20'b01010001110100010101: color_data = 12'b111011101110;
20'b01010001110100010110: color_data = 12'b111011101110;
20'b01010001110100010111: color_data = 12'b111011101110;
20'b01010001110100011001: color_data = 12'b111011101110;
20'b01010001110100011010: color_data = 12'b111011101110;
20'b01010001110100011011: color_data = 12'b111011101110;
20'b01010001110100011100: color_data = 12'b111011101110;
20'b01010001110100011101: color_data = 12'b111011101110;
20'b01010001110100011110: color_data = 12'b111011101110;
20'b01010001110100011111: color_data = 12'b111011101110;
20'b01010001110100100000: color_data = 12'b111011101110;
20'b01010001110100100001: color_data = 12'b111011101110;
20'b01010001110100100010: color_data = 12'b111011101110;
20'b01010001110100100100: color_data = 12'b111011101110;
20'b01010001110100100101: color_data = 12'b111011101110;
20'b01010001110100100110: color_data = 12'b111011101110;
20'b01010001110100100111: color_data = 12'b111011101110;
20'b01010001110100101000: color_data = 12'b111011101110;
20'b01010001110100101001: color_data = 12'b111011101110;
20'b01010001110100101010: color_data = 12'b111011101110;
20'b01010001110100101011: color_data = 12'b111011101110;
20'b01010001110100101100: color_data = 12'b111011101110;
20'b01010001110100101101: color_data = 12'b111011101110;
20'b01010001110101000100: color_data = 12'b111011101110;
20'b01010001110101000101: color_data = 12'b111011101110;
20'b01010001110101000110: color_data = 12'b111011101110;
20'b01010001110101000111: color_data = 12'b111011101110;
20'b01010001110101001000: color_data = 12'b111011101110;
20'b01010001110101001001: color_data = 12'b111011101110;
20'b01010001110101001010: color_data = 12'b111011101110;
20'b01010001110101001011: color_data = 12'b111011101110;
20'b01010001110101001100: color_data = 12'b111011101110;
20'b01010001110101001101: color_data = 12'b111011101110;
20'b01010001110101001111: color_data = 12'b111011101110;
20'b01010001110101010000: color_data = 12'b111011101110;
20'b01010001110101010001: color_data = 12'b111011101110;
20'b01010001110101010010: color_data = 12'b111011101110;
20'b01010001110101010011: color_data = 12'b111011101110;
20'b01010001110101010100: color_data = 12'b111011101110;
20'b01010001110101010101: color_data = 12'b111011101110;
20'b01010001110101010110: color_data = 12'b111011101110;
20'b01010001110101010111: color_data = 12'b111011101110;
20'b01010001110101011000: color_data = 12'b111011101110;
20'b01010001110101011010: color_data = 12'b111011101110;
20'b01010001110101011011: color_data = 12'b111011101110;
20'b01010001110101011100: color_data = 12'b111011101110;
20'b01010001110101011101: color_data = 12'b111011101110;
20'b01010001110101011110: color_data = 12'b111011101110;
20'b01010001110101011111: color_data = 12'b111011101110;
20'b01010001110101100000: color_data = 12'b111011101110;
20'b01010001110101100001: color_data = 12'b111011101110;
20'b01010001110101100010: color_data = 12'b111011101110;
20'b01010001110101100011: color_data = 12'b111011101110;
20'b01010001110101100101: color_data = 12'b111011101110;
20'b01010001110101100110: color_data = 12'b111011101110;
20'b01010001110101100111: color_data = 12'b111011101110;
20'b01010001110101101000: color_data = 12'b111011101110;
20'b01010001110101101001: color_data = 12'b111011101110;
20'b01010001110101101010: color_data = 12'b111011101110;
20'b01010001110101101011: color_data = 12'b111011101110;
20'b01010001110101101100: color_data = 12'b111011101110;
20'b01010001110101101101: color_data = 12'b111011101110;
20'b01010001110101101110: color_data = 12'b111011101110;
20'b01010001110101110000: color_data = 12'b111011101110;
20'b01010001110101110001: color_data = 12'b111011101110;
20'b01010001110101110010: color_data = 12'b111011101110;
20'b01010001110101110011: color_data = 12'b111011101110;
20'b01010001110101110100: color_data = 12'b111011101110;
20'b01010001110101110101: color_data = 12'b111011101110;
20'b01010001110101110110: color_data = 12'b111011101110;
20'b01010001110101110111: color_data = 12'b111011101110;
20'b01010001110101111000: color_data = 12'b111011101110;
20'b01010001110101111001: color_data = 12'b111011101110;
20'b01010001110101111011: color_data = 12'b111011101110;
20'b01010001110101111100: color_data = 12'b111011101110;
20'b01010001110101111101: color_data = 12'b111011101110;
20'b01010001110101111110: color_data = 12'b111011101110;
20'b01010001110101111111: color_data = 12'b111011101110;
20'b01010001110110000000: color_data = 12'b111011101110;
20'b01010001110110000001: color_data = 12'b111011101110;
20'b01010001110110000010: color_data = 12'b111011101110;
20'b01010001110110000011: color_data = 12'b111011101110;
20'b01010001110110000100: color_data = 12'b111011101110;
20'b01010001110110000110: color_data = 12'b111011101110;
20'b01010001110110000111: color_data = 12'b111011101110;
20'b01010001110110001000: color_data = 12'b111011101110;
20'b01010001110110001001: color_data = 12'b111011101110;
20'b01010001110110001010: color_data = 12'b111011101110;
20'b01010001110110001011: color_data = 12'b111011101110;
20'b01010001110110001100: color_data = 12'b111011101110;
20'b01010001110110001101: color_data = 12'b111011101110;
20'b01010001110110001110: color_data = 12'b111011101110;
20'b01010001110110001111: color_data = 12'b111011101110;
20'b01010001110110011100: color_data = 12'b111011101110;
20'b01010001110110011101: color_data = 12'b111011101110;
20'b01010001110110011110: color_data = 12'b111011101110;
20'b01010001110110011111: color_data = 12'b111011101110;
20'b01010001110110100000: color_data = 12'b111011101110;
20'b01010001110110100001: color_data = 12'b111011101110;
20'b01010001110110100010: color_data = 12'b111011101110;
20'b01010001110110100011: color_data = 12'b111011101110;
20'b01010001110110100100: color_data = 12'b111011101110;
20'b01010001110110100101: color_data = 12'b111011101110;
20'b01010001110110100111: color_data = 12'b111011101110;
20'b01010001110110101000: color_data = 12'b111011101110;
20'b01010001110110101001: color_data = 12'b111011101110;
20'b01010001110110101010: color_data = 12'b111011101110;
20'b01010001110110101011: color_data = 12'b111011101110;
20'b01010001110110101100: color_data = 12'b111011101110;
20'b01010001110110101101: color_data = 12'b111011101110;
20'b01010001110110101110: color_data = 12'b111011101110;
20'b01010001110110101111: color_data = 12'b111011101110;
20'b01010001110110110000: color_data = 12'b111011101110;
20'b01010001110111001000: color_data = 12'b111011101110;
20'b01010001110111001001: color_data = 12'b111011101110;
20'b01010001110111001010: color_data = 12'b111011101110;
20'b01010001110111001011: color_data = 12'b111011101110;
20'b01010001110111001100: color_data = 12'b111011101110;
20'b01010001110111001101: color_data = 12'b111011101110;
20'b01010001110111001110: color_data = 12'b111011101110;
20'b01010001110111001111: color_data = 12'b111011101110;
20'b01010001110111010000: color_data = 12'b111011101110;
20'b01010001110111010001: color_data = 12'b111011101110;
20'b01010001110111010011: color_data = 12'b111011101110;
20'b01010001110111010100: color_data = 12'b111011101110;
20'b01010001110111010101: color_data = 12'b111011101110;
20'b01010001110111010110: color_data = 12'b111011101110;
20'b01010001110111010111: color_data = 12'b111011101110;
20'b01010001110111011000: color_data = 12'b111011101110;
20'b01010001110111011001: color_data = 12'b111011101110;
20'b01010001110111011010: color_data = 12'b111011101110;
20'b01010001110111011011: color_data = 12'b111011101110;
20'b01010001110111011100: color_data = 12'b111011101110;
20'b01010010000010100001: color_data = 12'b111011101110;
20'b01010010000010100010: color_data = 12'b111011101110;
20'b01010010000010100011: color_data = 12'b111011101110;
20'b01010010000010100100: color_data = 12'b111011101110;
20'b01010010000010100101: color_data = 12'b111011101110;
20'b01010010000010100110: color_data = 12'b111011101110;
20'b01010010000010100111: color_data = 12'b111011101110;
20'b01010010000010101000: color_data = 12'b111011101110;
20'b01010010000010101001: color_data = 12'b111011101110;
20'b01010010000010101010: color_data = 12'b111011101110;
20'b01010010000010101100: color_data = 12'b111011101110;
20'b01010010000010101101: color_data = 12'b111011101110;
20'b01010010000010101110: color_data = 12'b111011101110;
20'b01010010000010101111: color_data = 12'b111011101110;
20'b01010010000010110000: color_data = 12'b111011101110;
20'b01010010000010110001: color_data = 12'b111011101110;
20'b01010010000010110010: color_data = 12'b111011101110;
20'b01010010000010110011: color_data = 12'b111011101110;
20'b01010010000010110100: color_data = 12'b111011101110;
20'b01010010000010110101: color_data = 12'b111011101110;
20'b01010010000010110111: color_data = 12'b111011101110;
20'b01010010000010111000: color_data = 12'b111011101110;
20'b01010010000010111001: color_data = 12'b111011101110;
20'b01010010000010111010: color_data = 12'b111011101110;
20'b01010010000010111011: color_data = 12'b111011101110;
20'b01010010000010111100: color_data = 12'b111011101110;
20'b01010010000010111101: color_data = 12'b111011101110;
20'b01010010000010111110: color_data = 12'b111011101110;
20'b01010010000010111111: color_data = 12'b111011101110;
20'b01010010000011000000: color_data = 12'b111011101110;
20'b01010010000011000010: color_data = 12'b111011101110;
20'b01010010000011000011: color_data = 12'b111011101110;
20'b01010010000011000100: color_data = 12'b111011101110;
20'b01010010000011000101: color_data = 12'b111011101110;
20'b01010010000011000110: color_data = 12'b111011101110;
20'b01010010000011000111: color_data = 12'b111011101110;
20'b01010010000011001000: color_data = 12'b111011101110;
20'b01010010000011001001: color_data = 12'b111011101110;
20'b01010010000011001010: color_data = 12'b111011101110;
20'b01010010000011001011: color_data = 12'b111011101110;
20'b01010010000011001101: color_data = 12'b111011101110;
20'b01010010000011001110: color_data = 12'b111011101110;
20'b01010010000011001111: color_data = 12'b111011101110;
20'b01010010000011010000: color_data = 12'b111011101110;
20'b01010010000011010001: color_data = 12'b111011101110;
20'b01010010000011010010: color_data = 12'b111011101110;
20'b01010010000011010011: color_data = 12'b111011101110;
20'b01010010000011010100: color_data = 12'b111011101110;
20'b01010010000011010101: color_data = 12'b111011101110;
20'b01010010000011010110: color_data = 12'b111011101110;
20'b01010010000011111000: color_data = 12'b111011101110;
20'b01010010000011111001: color_data = 12'b111011101110;
20'b01010010000011111010: color_data = 12'b111011101110;
20'b01010010000011111011: color_data = 12'b111011101110;
20'b01010010000011111100: color_data = 12'b111011101110;
20'b01010010000011111101: color_data = 12'b111011101110;
20'b01010010000011111110: color_data = 12'b111011101110;
20'b01010010000011111111: color_data = 12'b111011101110;
20'b01010010000100000000: color_data = 12'b111011101110;
20'b01010010000100000001: color_data = 12'b111011101110;
20'b01010010000100000011: color_data = 12'b111011101110;
20'b01010010000100000100: color_data = 12'b111011101110;
20'b01010010000100000101: color_data = 12'b111011101110;
20'b01010010000100000110: color_data = 12'b111011101110;
20'b01010010000100000111: color_data = 12'b111011101110;
20'b01010010000100001000: color_data = 12'b111011101110;
20'b01010010000100001001: color_data = 12'b111011101110;
20'b01010010000100001010: color_data = 12'b111011101110;
20'b01010010000100001011: color_data = 12'b111011101110;
20'b01010010000100001100: color_data = 12'b111011101110;
20'b01010010000100001110: color_data = 12'b111011101110;
20'b01010010000100001111: color_data = 12'b111011101110;
20'b01010010000100010000: color_data = 12'b111011101110;
20'b01010010000100010001: color_data = 12'b111011101110;
20'b01010010000100010010: color_data = 12'b111011101110;
20'b01010010000100010011: color_data = 12'b111011101110;
20'b01010010000100010100: color_data = 12'b111011101110;
20'b01010010000100010101: color_data = 12'b111011101110;
20'b01010010000100010110: color_data = 12'b111011101110;
20'b01010010000100010111: color_data = 12'b111011101110;
20'b01010010000100011001: color_data = 12'b111011101110;
20'b01010010000100011010: color_data = 12'b111011101110;
20'b01010010000100011011: color_data = 12'b111011101110;
20'b01010010000100011100: color_data = 12'b111011101110;
20'b01010010000100011101: color_data = 12'b111011101110;
20'b01010010000100011110: color_data = 12'b111011101110;
20'b01010010000100011111: color_data = 12'b111011101110;
20'b01010010000100100000: color_data = 12'b111011101110;
20'b01010010000100100001: color_data = 12'b111011101110;
20'b01010010000100100010: color_data = 12'b111011101110;
20'b01010010000100100100: color_data = 12'b111011101110;
20'b01010010000100100101: color_data = 12'b111011101110;
20'b01010010000100100110: color_data = 12'b111011101110;
20'b01010010000100100111: color_data = 12'b111011101110;
20'b01010010000100101000: color_data = 12'b111011101110;
20'b01010010000100101001: color_data = 12'b111011101110;
20'b01010010000100101010: color_data = 12'b111011101110;
20'b01010010000100101011: color_data = 12'b111011101110;
20'b01010010000100101100: color_data = 12'b111011101110;
20'b01010010000100101101: color_data = 12'b111011101110;
20'b01010010000101000100: color_data = 12'b111011101110;
20'b01010010000101000101: color_data = 12'b111011101110;
20'b01010010000101000110: color_data = 12'b111011101110;
20'b01010010000101000111: color_data = 12'b111011101110;
20'b01010010000101001000: color_data = 12'b111011101110;
20'b01010010000101001001: color_data = 12'b111011101110;
20'b01010010000101001010: color_data = 12'b111011101110;
20'b01010010000101001011: color_data = 12'b111011101110;
20'b01010010000101001100: color_data = 12'b111011101110;
20'b01010010000101001101: color_data = 12'b111011101110;
20'b01010010000101001111: color_data = 12'b111011101110;
20'b01010010000101010000: color_data = 12'b111011101110;
20'b01010010000101010001: color_data = 12'b111011101110;
20'b01010010000101010010: color_data = 12'b111011101110;
20'b01010010000101010011: color_data = 12'b111011101110;
20'b01010010000101010100: color_data = 12'b111011101110;
20'b01010010000101010101: color_data = 12'b111011101110;
20'b01010010000101010110: color_data = 12'b111011101110;
20'b01010010000101010111: color_data = 12'b111011101110;
20'b01010010000101011000: color_data = 12'b111011101110;
20'b01010010000101011010: color_data = 12'b111011101110;
20'b01010010000101011011: color_data = 12'b111011101110;
20'b01010010000101011100: color_data = 12'b111011101110;
20'b01010010000101011101: color_data = 12'b111011101110;
20'b01010010000101011110: color_data = 12'b111011101110;
20'b01010010000101011111: color_data = 12'b111011101110;
20'b01010010000101100000: color_data = 12'b111011101110;
20'b01010010000101100001: color_data = 12'b111011101110;
20'b01010010000101100010: color_data = 12'b111011101110;
20'b01010010000101100011: color_data = 12'b111011101110;
20'b01010010000101100101: color_data = 12'b111011101110;
20'b01010010000101100110: color_data = 12'b111011101110;
20'b01010010000101100111: color_data = 12'b111011101110;
20'b01010010000101101000: color_data = 12'b111011101110;
20'b01010010000101101001: color_data = 12'b111011101110;
20'b01010010000101101010: color_data = 12'b111011101110;
20'b01010010000101101011: color_data = 12'b111011101110;
20'b01010010000101101100: color_data = 12'b111011101110;
20'b01010010000101101101: color_data = 12'b111011101110;
20'b01010010000101101110: color_data = 12'b111011101110;
20'b01010010000101110000: color_data = 12'b111011101110;
20'b01010010000101110001: color_data = 12'b111011101110;
20'b01010010000101110010: color_data = 12'b111011101110;
20'b01010010000101110011: color_data = 12'b111011101110;
20'b01010010000101110100: color_data = 12'b111011101110;
20'b01010010000101110101: color_data = 12'b111011101110;
20'b01010010000101110110: color_data = 12'b111011101110;
20'b01010010000101110111: color_data = 12'b111011101110;
20'b01010010000101111000: color_data = 12'b111011101110;
20'b01010010000101111001: color_data = 12'b111011101110;
20'b01010010000101111011: color_data = 12'b111011101110;
20'b01010010000101111100: color_data = 12'b111011101110;
20'b01010010000101111101: color_data = 12'b111011101110;
20'b01010010000101111110: color_data = 12'b111011101110;
20'b01010010000101111111: color_data = 12'b111011101110;
20'b01010010000110000000: color_data = 12'b111011101110;
20'b01010010000110000001: color_data = 12'b111011101110;
20'b01010010000110000010: color_data = 12'b111011101110;
20'b01010010000110000011: color_data = 12'b111011101110;
20'b01010010000110000100: color_data = 12'b111011101110;
20'b01010010000110000110: color_data = 12'b111011101110;
20'b01010010000110000111: color_data = 12'b111011101110;
20'b01010010000110001000: color_data = 12'b111011101110;
20'b01010010000110001001: color_data = 12'b111011101110;
20'b01010010000110001010: color_data = 12'b111011101110;
20'b01010010000110001011: color_data = 12'b111011101110;
20'b01010010000110001100: color_data = 12'b111011101110;
20'b01010010000110001101: color_data = 12'b111011101110;
20'b01010010000110001110: color_data = 12'b111011101110;
20'b01010010000110001111: color_data = 12'b111011101110;
20'b01010010000110011100: color_data = 12'b111011101110;
20'b01010010000110011101: color_data = 12'b111011101110;
20'b01010010000110011110: color_data = 12'b111011101110;
20'b01010010000110011111: color_data = 12'b111011101110;
20'b01010010000110100000: color_data = 12'b111011101110;
20'b01010010000110100001: color_data = 12'b111011101110;
20'b01010010000110100010: color_data = 12'b111011101110;
20'b01010010000110100011: color_data = 12'b111011101110;
20'b01010010000110100100: color_data = 12'b111011101110;
20'b01010010000110100101: color_data = 12'b111011101110;
20'b01010010000110100111: color_data = 12'b111011101110;
20'b01010010000110101000: color_data = 12'b111011101110;
20'b01010010000110101001: color_data = 12'b111011101110;
20'b01010010000110101010: color_data = 12'b111011101110;
20'b01010010000110101011: color_data = 12'b111011101110;
20'b01010010000110101100: color_data = 12'b111011101110;
20'b01010010000110101101: color_data = 12'b111011101110;
20'b01010010000110101110: color_data = 12'b111011101110;
20'b01010010000110101111: color_data = 12'b111011101110;
20'b01010010000110110000: color_data = 12'b111011101110;
20'b01010010000111001000: color_data = 12'b111011101110;
20'b01010010000111001001: color_data = 12'b111011101110;
20'b01010010000111001010: color_data = 12'b111011101110;
20'b01010010000111001011: color_data = 12'b111011101110;
20'b01010010000111001100: color_data = 12'b111011101110;
20'b01010010000111001101: color_data = 12'b111011101110;
20'b01010010000111001110: color_data = 12'b111011101110;
20'b01010010000111001111: color_data = 12'b111011101110;
20'b01010010000111010000: color_data = 12'b111011101110;
20'b01010010000111010001: color_data = 12'b111011101110;
20'b01010010000111010011: color_data = 12'b111011101110;
20'b01010010000111010100: color_data = 12'b111011101110;
20'b01010010000111010101: color_data = 12'b111011101110;
20'b01010010000111010110: color_data = 12'b111011101110;
20'b01010010000111010111: color_data = 12'b111011101110;
20'b01010010000111011000: color_data = 12'b111011101110;
20'b01010010000111011001: color_data = 12'b111011101110;
20'b01010010000111011010: color_data = 12'b111011101110;
20'b01010010000111011011: color_data = 12'b111011101110;
20'b01010010000111011100: color_data = 12'b111011101110;
20'b01010010010010100001: color_data = 12'b111011101110;
20'b01010010010010100010: color_data = 12'b111011101110;
20'b01010010010010100011: color_data = 12'b111011101110;
20'b01010010010010100100: color_data = 12'b111011101110;
20'b01010010010010100101: color_data = 12'b111011101110;
20'b01010010010010100110: color_data = 12'b111011101110;
20'b01010010010010100111: color_data = 12'b111011101110;
20'b01010010010010101000: color_data = 12'b111011101110;
20'b01010010010010101001: color_data = 12'b111011101110;
20'b01010010010010101010: color_data = 12'b111011101110;
20'b01010010010010101100: color_data = 12'b111011101110;
20'b01010010010010101101: color_data = 12'b111011101110;
20'b01010010010010101110: color_data = 12'b111011101110;
20'b01010010010010101111: color_data = 12'b111011101110;
20'b01010010010010110000: color_data = 12'b111011101110;
20'b01010010010010110001: color_data = 12'b111011101110;
20'b01010010010010110010: color_data = 12'b111011101110;
20'b01010010010010110011: color_data = 12'b111011101110;
20'b01010010010010110100: color_data = 12'b111011101110;
20'b01010010010010110101: color_data = 12'b111011101110;
20'b01010010010010110111: color_data = 12'b111011101110;
20'b01010010010010111000: color_data = 12'b111011101110;
20'b01010010010010111001: color_data = 12'b111011101110;
20'b01010010010010111010: color_data = 12'b111011101110;
20'b01010010010010111011: color_data = 12'b111011101110;
20'b01010010010010111100: color_data = 12'b111011101110;
20'b01010010010010111101: color_data = 12'b111011101110;
20'b01010010010010111110: color_data = 12'b111011101110;
20'b01010010010010111111: color_data = 12'b111011101110;
20'b01010010010011000000: color_data = 12'b111011101110;
20'b01010010010011000010: color_data = 12'b111011101110;
20'b01010010010011000011: color_data = 12'b111011101110;
20'b01010010010011000100: color_data = 12'b111011101110;
20'b01010010010011000101: color_data = 12'b111011101110;
20'b01010010010011000110: color_data = 12'b111011101110;
20'b01010010010011000111: color_data = 12'b111011101110;
20'b01010010010011001000: color_data = 12'b111011101110;
20'b01010010010011001001: color_data = 12'b111011101110;
20'b01010010010011001010: color_data = 12'b111011101110;
20'b01010010010011001011: color_data = 12'b111011101110;
20'b01010010010011001101: color_data = 12'b111011101110;
20'b01010010010011001110: color_data = 12'b111011101110;
20'b01010010010011001111: color_data = 12'b111011101110;
20'b01010010010011010000: color_data = 12'b111011101110;
20'b01010010010011010001: color_data = 12'b111011101110;
20'b01010010010011010010: color_data = 12'b111011101110;
20'b01010010010011010011: color_data = 12'b111011101110;
20'b01010010010011010100: color_data = 12'b111011101110;
20'b01010010010011010101: color_data = 12'b111011101110;
20'b01010010010011010110: color_data = 12'b111011101110;
20'b01010010010011111000: color_data = 12'b111011101110;
20'b01010010010011111001: color_data = 12'b111011101110;
20'b01010010010011111010: color_data = 12'b111011101110;
20'b01010010010011111011: color_data = 12'b111011101110;
20'b01010010010011111100: color_data = 12'b111011101110;
20'b01010010010011111101: color_data = 12'b111011101110;
20'b01010010010011111110: color_data = 12'b111011101110;
20'b01010010010011111111: color_data = 12'b111011101110;
20'b01010010010100000000: color_data = 12'b111011101110;
20'b01010010010100000001: color_data = 12'b111011101110;
20'b01010010010100000011: color_data = 12'b111011101110;
20'b01010010010100000100: color_data = 12'b111011101110;
20'b01010010010100000101: color_data = 12'b111011101110;
20'b01010010010100000110: color_data = 12'b111011101110;
20'b01010010010100000111: color_data = 12'b111011101110;
20'b01010010010100001000: color_data = 12'b111011101110;
20'b01010010010100001001: color_data = 12'b111011101110;
20'b01010010010100001010: color_data = 12'b111011101110;
20'b01010010010100001011: color_data = 12'b111011101110;
20'b01010010010100001100: color_data = 12'b111011101110;
20'b01010010010100001110: color_data = 12'b111011101110;
20'b01010010010100001111: color_data = 12'b111011101110;
20'b01010010010100010000: color_data = 12'b111011101110;
20'b01010010010100010001: color_data = 12'b111011101110;
20'b01010010010100010010: color_data = 12'b111011101110;
20'b01010010010100010011: color_data = 12'b111011101110;
20'b01010010010100010100: color_data = 12'b111011101110;
20'b01010010010100010101: color_data = 12'b111011101110;
20'b01010010010100010110: color_data = 12'b111011101110;
20'b01010010010100010111: color_data = 12'b111011101110;
20'b01010010010100011001: color_data = 12'b111011101110;
20'b01010010010100011010: color_data = 12'b111011101110;
20'b01010010010100011011: color_data = 12'b111011101110;
20'b01010010010100011100: color_data = 12'b111011101110;
20'b01010010010100011101: color_data = 12'b111011101110;
20'b01010010010100011110: color_data = 12'b111011101110;
20'b01010010010100011111: color_data = 12'b111011101110;
20'b01010010010100100000: color_data = 12'b111011101110;
20'b01010010010100100001: color_data = 12'b111011101110;
20'b01010010010100100010: color_data = 12'b111011101110;
20'b01010010010100100100: color_data = 12'b111011101110;
20'b01010010010100100101: color_data = 12'b111011101110;
20'b01010010010100100110: color_data = 12'b111011101110;
20'b01010010010100100111: color_data = 12'b111011101110;
20'b01010010010100101000: color_data = 12'b111011101110;
20'b01010010010100101001: color_data = 12'b111011101110;
20'b01010010010100101010: color_data = 12'b111011101110;
20'b01010010010100101011: color_data = 12'b111011101110;
20'b01010010010100101100: color_data = 12'b111011101110;
20'b01010010010100101101: color_data = 12'b111011101110;
20'b01010010010101000100: color_data = 12'b111011101110;
20'b01010010010101000101: color_data = 12'b111011101110;
20'b01010010010101000110: color_data = 12'b111011101110;
20'b01010010010101000111: color_data = 12'b111011101110;
20'b01010010010101001000: color_data = 12'b111011101110;
20'b01010010010101001001: color_data = 12'b111011101110;
20'b01010010010101001010: color_data = 12'b111011101110;
20'b01010010010101001011: color_data = 12'b111011101110;
20'b01010010010101001100: color_data = 12'b111011101110;
20'b01010010010101001101: color_data = 12'b111011101110;
20'b01010010010101001111: color_data = 12'b111011101110;
20'b01010010010101010000: color_data = 12'b111011101110;
20'b01010010010101010001: color_data = 12'b111011101110;
20'b01010010010101010010: color_data = 12'b111011101110;
20'b01010010010101010011: color_data = 12'b111011101110;
20'b01010010010101010100: color_data = 12'b111011101110;
20'b01010010010101010101: color_data = 12'b111011101110;
20'b01010010010101010110: color_data = 12'b111011101110;
20'b01010010010101010111: color_data = 12'b111011101110;
20'b01010010010101011000: color_data = 12'b111011101110;
20'b01010010010101011010: color_data = 12'b111011101110;
20'b01010010010101011011: color_data = 12'b111011101110;
20'b01010010010101011100: color_data = 12'b111011101110;
20'b01010010010101011101: color_data = 12'b111011101110;
20'b01010010010101011110: color_data = 12'b111011101110;
20'b01010010010101011111: color_data = 12'b111011101110;
20'b01010010010101100000: color_data = 12'b111011101110;
20'b01010010010101100001: color_data = 12'b111011101110;
20'b01010010010101100010: color_data = 12'b111011101110;
20'b01010010010101100011: color_data = 12'b111011101110;
20'b01010010010101100101: color_data = 12'b111011101110;
20'b01010010010101100110: color_data = 12'b111011101110;
20'b01010010010101100111: color_data = 12'b111011101110;
20'b01010010010101101000: color_data = 12'b111011101110;
20'b01010010010101101001: color_data = 12'b111011101110;
20'b01010010010101101010: color_data = 12'b111011101110;
20'b01010010010101101011: color_data = 12'b111011101110;
20'b01010010010101101100: color_data = 12'b111011101110;
20'b01010010010101101101: color_data = 12'b111011101110;
20'b01010010010101101110: color_data = 12'b111011101110;
20'b01010010010101110000: color_data = 12'b111011101110;
20'b01010010010101110001: color_data = 12'b111011101110;
20'b01010010010101110010: color_data = 12'b111011101110;
20'b01010010010101110011: color_data = 12'b111011101110;
20'b01010010010101110100: color_data = 12'b111011101110;
20'b01010010010101110101: color_data = 12'b111011101110;
20'b01010010010101110110: color_data = 12'b111011101110;
20'b01010010010101110111: color_data = 12'b111011101110;
20'b01010010010101111000: color_data = 12'b111011101110;
20'b01010010010101111001: color_data = 12'b111011101110;
20'b01010010010101111011: color_data = 12'b111011101110;
20'b01010010010101111100: color_data = 12'b111011101110;
20'b01010010010101111101: color_data = 12'b111011101110;
20'b01010010010101111110: color_data = 12'b111011101110;
20'b01010010010101111111: color_data = 12'b111011101110;
20'b01010010010110000000: color_data = 12'b111011101110;
20'b01010010010110000001: color_data = 12'b111011101110;
20'b01010010010110000010: color_data = 12'b111011101110;
20'b01010010010110000011: color_data = 12'b111011101110;
20'b01010010010110000100: color_data = 12'b111011101110;
20'b01010010010110000110: color_data = 12'b111011101110;
20'b01010010010110000111: color_data = 12'b111011101110;
20'b01010010010110001000: color_data = 12'b111011101110;
20'b01010010010110001001: color_data = 12'b111011101110;
20'b01010010010110001010: color_data = 12'b111011101110;
20'b01010010010110001011: color_data = 12'b111011101110;
20'b01010010010110001100: color_data = 12'b111011101110;
20'b01010010010110001101: color_data = 12'b111011101110;
20'b01010010010110001110: color_data = 12'b111011101110;
20'b01010010010110001111: color_data = 12'b111011101110;
20'b01010010010110011100: color_data = 12'b111011101110;
20'b01010010010110011101: color_data = 12'b111011101110;
20'b01010010010110011110: color_data = 12'b111011101110;
20'b01010010010110011111: color_data = 12'b111011101110;
20'b01010010010110100000: color_data = 12'b111011101110;
20'b01010010010110100001: color_data = 12'b111011101110;
20'b01010010010110100010: color_data = 12'b111011101110;
20'b01010010010110100011: color_data = 12'b111011101110;
20'b01010010010110100100: color_data = 12'b111011101110;
20'b01010010010110100101: color_data = 12'b111011101110;
20'b01010010010110100111: color_data = 12'b111011101110;
20'b01010010010110101000: color_data = 12'b111011101110;
20'b01010010010110101001: color_data = 12'b111011101110;
20'b01010010010110101010: color_data = 12'b111011101110;
20'b01010010010110101011: color_data = 12'b111011101110;
20'b01010010010110101100: color_data = 12'b111011101110;
20'b01010010010110101101: color_data = 12'b111011101110;
20'b01010010010110101110: color_data = 12'b111011101110;
20'b01010010010110101111: color_data = 12'b111011101110;
20'b01010010010110110000: color_data = 12'b111011101110;
20'b01010010010111001000: color_data = 12'b111011101110;
20'b01010010010111001001: color_data = 12'b111011101110;
20'b01010010010111001010: color_data = 12'b111011101110;
20'b01010010010111001011: color_data = 12'b111011101110;
20'b01010010010111001100: color_data = 12'b111011101110;
20'b01010010010111001101: color_data = 12'b111011101110;
20'b01010010010111001110: color_data = 12'b111011101110;
20'b01010010010111001111: color_data = 12'b111011101110;
20'b01010010010111010000: color_data = 12'b111011101110;
20'b01010010010111010001: color_data = 12'b111011101110;
20'b01010010010111010011: color_data = 12'b111011101110;
20'b01010010010111010100: color_data = 12'b111011101110;
20'b01010010010111010101: color_data = 12'b111011101110;
20'b01010010010111010110: color_data = 12'b111011101110;
20'b01010010010111010111: color_data = 12'b111011101110;
20'b01010010010111011000: color_data = 12'b111011101110;
20'b01010010010111011001: color_data = 12'b111011101110;
20'b01010010010111011010: color_data = 12'b111011101110;
20'b01010010010111011011: color_data = 12'b111011101110;
20'b01010010010111011100: color_data = 12'b111011101110;
20'b01010010100010100001: color_data = 12'b111011101110;
20'b01010010100010100010: color_data = 12'b111011101110;
20'b01010010100010100011: color_data = 12'b111011101110;
20'b01010010100010100100: color_data = 12'b111011101110;
20'b01010010100010100101: color_data = 12'b111011101110;
20'b01010010100010100110: color_data = 12'b111011101110;
20'b01010010100010100111: color_data = 12'b111011101110;
20'b01010010100010101000: color_data = 12'b111011101110;
20'b01010010100010101001: color_data = 12'b111011101110;
20'b01010010100010101010: color_data = 12'b111011101110;
20'b01010010100010101100: color_data = 12'b111011101110;
20'b01010010100010101101: color_data = 12'b111011101110;
20'b01010010100010101110: color_data = 12'b111011101110;
20'b01010010100010101111: color_data = 12'b111011101110;
20'b01010010100010110000: color_data = 12'b111011101110;
20'b01010010100010110001: color_data = 12'b111011101110;
20'b01010010100010110010: color_data = 12'b111011101110;
20'b01010010100010110011: color_data = 12'b111011101110;
20'b01010010100010110100: color_data = 12'b111011101110;
20'b01010010100010110101: color_data = 12'b111011101110;
20'b01010010100010110111: color_data = 12'b111011101110;
20'b01010010100010111000: color_data = 12'b111011101110;
20'b01010010100010111001: color_data = 12'b111011101110;
20'b01010010100010111010: color_data = 12'b111011101110;
20'b01010010100010111011: color_data = 12'b111011101110;
20'b01010010100010111100: color_data = 12'b111011101110;
20'b01010010100010111101: color_data = 12'b111011101110;
20'b01010010100010111110: color_data = 12'b111011101110;
20'b01010010100010111111: color_data = 12'b111011101110;
20'b01010010100011000000: color_data = 12'b111011101110;
20'b01010010100011000010: color_data = 12'b111011101110;
20'b01010010100011000011: color_data = 12'b111011101110;
20'b01010010100011000100: color_data = 12'b111011101110;
20'b01010010100011000101: color_data = 12'b111011101110;
20'b01010010100011000110: color_data = 12'b111011101110;
20'b01010010100011000111: color_data = 12'b111011101110;
20'b01010010100011001000: color_data = 12'b111011101110;
20'b01010010100011001001: color_data = 12'b111011101110;
20'b01010010100011001010: color_data = 12'b111011101110;
20'b01010010100011001011: color_data = 12'b111011101110;
20'b01010010100011001101: color_data = 12'b111011101110;
20'b01010010100011001110: color_data = 12'b111011101110;
20'b01010010100011001111: color_data = 12'b111011101110;
20'b01010010100011010000: color_data = 12'b111011101110;
20'b01010010100011010001: color_data = 12'b111011101110;
20'b01010010100011010010: color_data = 12'b111011101110;
20'b01010010100011010011: color_data = 12'b111011101110;
20'b01010010100011010100: color_data = 12'b111011101110;
20'b01010010100011010101: color_data = 12'b111011101110;
20'b01010010100011010110: color_data = 12'b111011101110;
20'b01010010100011111000: color_data = 12'b111011101110;
20'b01010010100011111001: color_data = 12'b111011101110;
20'b01010010100011111010: color_data = 12'b111011101110;
20'b01010010100011111011: color_data = 12'b111011101110;
20'b01010010100011111100: color_data = 12'b111011101110;
20'b01010010100011111101: color_data = 12'b111011101110;
20'b01010010100011111110: color_data = 12'b111011101110;
20'b01010010100011111111: color_data = 12'b111011101110;
20'b01010010100100000000: color_data = 12'b111011101110;
20'b01010010100100000001: color_data = 12'b111011101110;
20'b01010010100100000011: color_data = 12'b111011101110;
20'b01010010100100000100: color_data = 12'b111011101110;
20'b01010010100100000101: color_data = 12'b111011101110;
20'b01010010100100000110: color_data = 12'b111011101110;
20'b01010010100100000111: color_data = 12'b111011101110;
20'b01010010100100001000: color_data = 12'b111011101110;
20'b01010010100100001001: color_data = 12'b111011101110;
20'b01010010100100001010: color_data = 12'b111011101110;
20'b01010010100100001011: color_data = 12'b111011101110;
20'b01010010100100001100: color_data = 12'b111011101110;
20'b01010010100100001110: color_data = 12'b111011101110;
20'b01010010100100001111: color_data = 12'b111011101110;
20'b01010010100100010000: color_data = 12'b111011101110;
20'b01010010100100010001: color_data = 12'b111011101110;
20'b01010010100100010010: color_data = 12'b111011101110;
20'b01010010100100010011: color_data = 12'b111011101110;
20'b01010010100100010100: color_data = 12'b111011101110;
20'b01010010100100010101: color_data = 12'b111011101110;
20'b01010010100100010110: color_data = 12'b111011101110;
20'b01010010100100010111: color_data = 12'b111011101110;
20'b01010010100100011001: color_data = 12'b111011101110;
20'b01010010100100011010: color_data = 12'b111011101110;
20'b01010010100100011011: color_data = 12'b111011101110;
20'b01010010100100011100: color_data = 12'b111011101110;
20'b01010010100100011101: color_data = 12'b111011101110;
20'b01010010100100011110: color_data = 12'b111011101110;
20'b01010010100100011111: color_data = 12'b111011101110;
20'b01010010100100100000: color_data = 12'b111011101110;
20'b01010010100100100001: color_data = 12'b111011101110;
20'b01010010100100100010: color_data = 12'b111011101110;
20'b01010010100100100100: color_data = 12'b111011101110;
20'b01010010100100100101: color_data = 12'b111011101110;
20'b01010010100100100110: color_data = 12'b111011101110;
20'b01010010100100100111: color_data = 12'b111011101110;
20'b01010010100100101000: color_data = 12'b111011101110;
20'b01010010100100101001: color_data = 12'b111011101110;
20'b01010010100100101010: color_data = 12'b111011101110;
20'b01010010100100101011: color_data = 12'b111011101110;
20'b01010010100100101100: color_data = 12'b111011101110;
20'b01010010100100101101: color_data = 12'b111011101110;
20'b01010010100101000100: color_data = 12'b111011101110;
20'b01010010100101000101: color_data = 12'b111011101110;
20'b01010010100101000110: color_data = 12'b111011101110;
20'b01010010100101000111: color_data = 12'b111011101110;
20'b01010010100101001000: color_data = 12'b111011101110;
20'b01010010100101001001: color_data = 12'b111011101110;
20'b01010010100101001010: color_data = 12'b111011101110;
20'b01010010100101001011: color_data = 12'b111011101110;
20'b01010010100101001100: color_data = 12'b111011101110;
20'b01010010100101001101: color_data = 12'b111011101110;
20'b01010010100101001111: color_data = 12'b111011101110;
20'b01010010100101010000: color_data = 12'b111011101110;
20'b01010010100101010001: color_data = 12'b111011101110;
20'b01010010100101010010: color_data = 12'b111011101110;
20'b01010010100101010011: color_data = 12'b111011101110;
20'b01010010100101010100: color_data = 12'b111011101110;
20'b01010010100101010101: color_data = 12'b111011101110;
20'b01010010100101010110: color_data = 12'b111011101110;
20'b01010010100101010111: color_data = 12'b111011101110;
20'b01010010100101011000: color_data = 12'b111011101110;
20'b01010010100101011010: color_data = 12'b111011101110;
20'b01010010100101011011: color_data = 12'b111011101110;
20'b01010010100101011100: color_data = 12'b111011101110;
20'b01010010100101011101: color_data = 12'b111011101110;
20'b01010010100101011110: color_data = 12'b111011101110;
20'b01010010100101011111: color_data = 12'b111011101110;
20'b01010010100101100000: color_data = 12'b111011101110;
20'b01010010100101100001: color_data = 12'b111011101110;
20'b01010010100101100010: color_data = 12'b111011101110;
20'b01010010100101100011: color_data = 12'b111011101110;
20'b01010010100101100101: color_data = 12'b111011101110;
20'b01010010100101100110: color_data = 12'b111011101110;
20'b01010010100101100111: color_data = 12'b111011101110;
20'b01010010100101101000: color_data = 12'b111011101110;
20'b01010010100101101001: color_data = 12'b111011101110;
20'b01010010100101101010: color_data = 12'b111011101110;
20'b01010010100101101011: color_data = 12'b111011101110;
20'b01010010100101101100: color_data = 12'b111011101110;
20'b01010010100101101101: color_data = 12'b111011101110;
20'b01010010100101101110: color_data = 12'b111011101110;
20'b01010010100101110000: color_data = 12'b111011101110;
20'b01010010100101110001: color_data = 12'b111011101110;
20'b01010010100101110010: color_data = 12'b111011101110;
20'b01010010100101110011: color_data = 12'b111011101110;
20'b01010010100101110100: color_data = 12'b111011101110;
20'b01010010100101110101: color_data = 12'b111011101110;
20'b01010010100101110110: color_data = 12'b111011101110;
20'b01010010100101110111: color_data = 12'b111011101110;
20'b01010010100101111000: color_data = 12'b111011101110;
20'b01010010100101111001: color_data = 12'b111011101110;
20'b01010010100101111011: color_data = 12'b111011101110;
20'b01010010100101111100: color_data = 12'b111011101110;
20'b01010010100101111101: color_data = 12'b111011101110;
20'b01010010100101111110: color_data = 12'b111011101110;
20'b01010010100101111111: color_data = 12'b111011101110;
20'b01010010100110000000: color_data = 12'b111011101110;
20'b01010010100110000001: color_data = 12'b111011101110;
20'b01010010100110000010: color_data = 12'b111011101110;
20'b01010010100110000011: color_data = 12'b111011101110;
20'b01010010100110000100: color_data = 12'b111011101110;
20'b01010010100110000110: color_data = 12'b111011101110;
20'b01010010100110000111: color_data = 12'b111011101110;
20'b01010010100110001000: color_data = 12'b111011101110;
20'b01010010100110001001: color_data = 12'b111011101110;
20'b01010010100110001010: color_data = 12'b111011101110;
20'b01010010100110001011: color_data = 12'b111011101110;
20'b01010010100110001100: color_data = 12'b111011101110;
20'b01010010100110001101: color_data = 12'b111011101110;
20'b01010010100110001110: color_data = 12'b111011101110;
20'b01010010100110001111: color_data = 12'b111011101110;
20'b01010010100110011100: color_data = 12'b111011101110;
20'b01010010100110011101: color_data = 12'b111011101110;
20'b01010010100110011110: color_data = 12'b111011101110;
20'b01010010100110011111: color_data = 12'b111011101110;
20'b01010010100110100000: color_data = 12'b111011101110;
20'b01010010100110100001: color_data = 12'b111011101110;
20'b01010010100110100010: color_data = 12'b111011101110;
20'b01010010100110100011: color_data = 12'b111011101110;
20'b01010010100110100100: color_data = 12'b111011101110;
20'b01010010100110100101: color_data = 12'b111011101110;
20'b01010010100110100111: color_data = 12'b111011101110;
20'b01010010100110101000: color_data = 12'b111011101110;
20'b01010010100110101001: color_data = 12'b111011101110;
20'b01010010100110101010: color_data = 12'b111011101110;
20'b01010010100110101011: color_data = 12'b111011101110;
20'b01010010100110101100: color_data = 12'b111011101110;
20'b01010010100110101101: color_data = 12'b111011101110;
20'b01010010100110101110: color_data = 12'b111011101110;
20'b01010010100110101111: color_data = 12'b111011101110;
20'b01010010100110110000: color_data = 12'b111011101110;
20'b01010010100111001000: color_data = 12'b111011101110;
20'b01010010100111001001: color_data = 12'b111011101110;
20'b01010010100111001010: color_data = 12'b111011101110;
20'b01010010100111001011: color_data = 12'b111011101110;
20'b01010010100111001100: color_data = 12'b111011101110;
20'b01010010100111001101: color_data = 12'b111011101110;
20'b01010010100111001110: color_data = 12'b111011101110;
20'b01010010100111001111: color_data = 12'b111011101110;
20'b01010010100111010000: color_data = 12'b111011101110;
20'b01010010100111010001: color_data = 12'b111011101110;
20'b01010010100111010011: color_data = 12'b111011101110;
20'b01010010100111010100: color_data = 12'b111011101110;
20'b01010010100111010101: color_data = 12'b111011101110;
20'b01010010100111010110: color_data = 12'b111011101110;
20'b01010010100111010111: color_data = 12'b111011101110;
20'b01010010100111011000: color_data = 12'b111011101110;
20'b01010010100111011001: color_data = 12'b111011101110;
20'b01010010100111011010: color_data = 12'b111011101110;
20'b01010010100111011011: color_data = 12'b111011101110;
20'b01010010100111011100: color_data = 12'b111011101110;
20'b01010010110010100001: color_data = 12'b111011101110;
20'b01010010110010100010: color_data = 12'b111011101110;
20'b01010010110010100011: color_data = 12'b111011101110;
20'b01010010110010100100: color_data = 12'b111011101110;
20'b01010010110010100101: color_data = 12'b111011101110;
20'b01010010110010100110: color_data = 12'b111011101110;
20'b01010010110010100111: color_data = 12'b111011101110;
20'b01010010110010101000: color_data = 12'b111011101110;
20'b01010010110010101001: color_data = 12'b111011101110;
20'b01010010110010101010: color_data = 12'b111011101110;
20'b01010010110010101100: color_data = 12'b111011101110;
20'b01010010110010101101: color_data = 12'b111011101110;
20'b01010010110010101110: color_data = 12'b111011101110;
20'b01010010110010101111: color_data = 12'b111011101110;
20'b01010010110010110000: color_data = 12'b111011101110;
20'b01010010110010110001: color_data = 12'b111011101110;
20'b01010010110010110010: color_data = 12'b111011101110;
20'b01010010110010110011: color_data = 12'b111011101110;
20'b01010010110010110100: color_data = 12'b111011101110;
20'b01010010110010110101: color_data = 12'b111011101110;
20'b01010010110010110111: color_data = 12'b111011101110;
20'b01010010110010111000: color_data = 12'b111011101110;
20'b01010010110010111001: color_data = 12'b111011101110;
20'b01010010110010111010: color_data = 12'b111011101110;
20'b01010010110010111011: color_data = 12'b111011101110;
20'b01010010110010111100: color_data = 12'b111011101110;
20'b01010010110010111101: color_data = 12'b111011101110;
20'b01010010110010111110: color_data = 12'b111011101110;
20'b01010010110010111111: color_data = 12'b111011101110;
20'b01010010110011000000: color_data = 12'b111011101110;
20'b01010010110011000010: color_data = 12'b111011101110;
20'b01010010110011000011: color_data = 12'b111011101110;
20'b01010010110011000100: color_data = 12'b111011101110;
20'b01010010110011000101: color_data = 12'b111011101110;
20'b01010010110011000110: color_data = 12'b111011101110;
20'b01010010110011000111: color_data = 12'b111011101110;
20'b01010010110011001000: color_data = 12'b111011101110;
20'b01010010110011001001: color_data = 12'b111011101110;
20'b01010010110011001010: color_data = 12'b111011101110;
20'b01010010110011001011: color_data = 12'b111011101110;
20'b01010010110011001101: color_data = 12'b111011101110;
20'b01010010110011001110: color_data = 12'b111011101110;
20'b01010010110011001111: color_data = 12'b111011101110;
20'b01010010110011010000: color_data = 12'b111011101110;
20'b01010010110011010001: color_data = 12'b111011101110;
20'b01010010110011010010: color_data = 12'b111011101110;
20'b01010010110011010011: color_data = 12'b111011101110;
20'b01010010110011010100: color_data = 12'b111011101110;
20'b01010010110011010101: color_data = 12'b111011101110;
20'b01010010110011010110: color_data = 12'b111011101110;
20'b01010010110011111000: color_data = 12'b111011101110;
20'b01010010110011111001: color_data = 12'b111011101110;
20'b01010010110011111010: color_data = 12'b111011101110;
20'b01010010110011111011: color_data = 12'b111011101110;
20'b01010010110011111100: color_data = 12'b111011101110;
20'b01010010110011111101: color_data = 12'b111011101110;
20'b01010010110011111110: color_data = 12'b111011101110;
20'b01010010110011111111: color_data = 12'b111011101110;
20'b01010010110100000000: color_data = 12'b111011101110;
20'b01010010110100000001: color_data = 12'b111011101110;
20'b01010010110100000011: color_data = 12'b111011101110;
20'b01010010110100000100: color_data = 12'b111011101110;
20'b01010010110100000101: color_data = 12'b111011101110;
20'b01010010110100000110: color_data = 12'b111011101110;
20'b01010010110100000111: color_data = 12'b111011101110;
20'b01010010110100001000: color_data = 12'b111011101110;
20'b01010010110100001001: color_data = 12'b111011101110;
20'b01010010110100001010: color_data = 12'b111011101110;
20'b01010010110100001011: color_data = 12'b111011101110;
20'b01010010110100001100: color_data = 12'b111011101110;
20'b01010010110100001110: color_data = 12'b111011101110;
20'b01010010110100001111: color_data = 12'b111011101110;
20'b01010010110100010000: color_data = 12'b111011101110;
20'b01010010110100010001: color_data = 12'b111011101110;
20'b01010010110100010010: color_data = 12'b111011101110;
20'b01010010110100010011: color_data = 12'b111011101110;
20'b01010010110100010100: color_data = 12'b111011101110;
20'b01010010110100010101: color_data = 12'b111011101110;
20'b01010010110100010110: color_data = 12'b111011101110;
20'b01010010110100010111: color_data = 12'b111011101110;
20'b01010010110100011001: color_data = 12'b111011101110;
20'b01010010110100011010: color_data = 12'b111011101110;
20'b01010010110100011011: color_data = 12'b111011101110;
20'b01010010110100011100: color_data = 12'b111011101110;
20'b01010010110100011101: color_data = 12'b111011101110;
20'b01010010110100011110: color_data = 12'b111011101110;
20'b01010010110100011111: color_data = 12'b111011101110;
20'b01010010110100100000: color_data = 12'b111011101110;
20'b01010010110100100001: color_data = 12'b111011101110;
20'b01010010110100100010: color_data = 12'b111011101110;
20'b01010010110100100100: color_data = 12'b111011101110;
20'b01010010110100100101: color_data = 12'b111011101110;
20'b01010010110100100110: color_data = 12'b111011101110;
20'b01010010110100100111: color_data = 12'b111011101110;
20'b01010010110100101000: color_data = 12'b111011101110;
20'b01010010110100101001: color_data = 12'b111011101110;
20'b01010010110100101010: color_data = 12'b111011101110;
20'b01010010110100101011: color_data = 12'b111011101110;
20'b01010010110100101100: color_data = 12'b111011101110;
20'b01010010110100101101: color_data = 12'b111011101110;
20'b01010010110101000100: color_data = 12'b111011101110;
20'b01010010110101000101: color_data = 12'b111011101110;
20'b01010010110101000110: color_data = 12'b111011101110;
20'b01010010110101000111: color_data = 12'b111011101110;
20'b01010010110101001000: color_data = 12'b111011101110;
20'b01010010110101001001: color_data = 12'b111011101110;
20'b01010010110101001010: color_data = 12'b111011101110;
20'b01010010110101001011: color_data = 12'b111011101110;
20'b01010010110101001100: color_data = 12'b111011101110;
20'b01010010110101001101: color_data = 12'b111011101110;
20'b01010010110101001111: color_data = 12'b111011101110;
20'b01010010110101010000: color_data = 12'b111011101110;
20'b01010010110101010001: color_data = 12'b111011101110;
20'b01010010110101010010: color_data = 12'b111011101110;
20'b01010010110101010011: color_data = 12'b111011101110;
20'b01010010110101010100: color_data = 12'b111011101110;
20'b01010010110101010101: color_data = 12'b111011101110;
20'b01010010110101010110: color_data = 12'b111011101110;
20'b01010010110101010111: color_data = 12'b111011101110;
20'b01010010110101011000: color_data = 12'b111011101110;
20'b01010010110101011010: color_data = 12'b111011101110;
20'b01010010110101011011: color_data = 12'b111011101110;
20'b01010010110101011100: color_data = 12'b111011101110;
20'b01010010110101011101: color_data = 12'b111011101110;
20'b01010010110101011110: color_data = 12'b111011101110;
20'b01010010110101011111: color_data = 12'b111011101110;
20'b01010010110101100000: color_data = 12'b111011101110;
20'b01010010110101100001: color_data = 12'b111011101110;
20'b01010010110101100010: color_data = 12'b111011101110;
20'b01010010110101100011: color_data = 12'b111011101110;
20'b01010010110101100101: color_data = 12'b111011101110;
20'b01010010110101100110: color_data = 12'b111011101110;
20'b01010010110101100111: color_data = 12'b111011101110;
20'b01010010110101101000: color_data = 12'b111011101110;
20'b01010010110101101001: color_data = 12'b111011101110;
20'b01010010110101101010: color_data = 12'b111011101110;
20'b01010010110101101011: color_data = 12'b111011101110;
20'b01010010110101101100: color_data = 12'b111011101110;
20'b01010010110101101101: color_data = 12'b111011101110;
20'b01010010110101101110: color_data = 12'b111011101110;
20'b01010010110101110000: color_data = 12'b111011101110;
20'b01010010110101110001: color_data = 12'b111011101110;
20'b01010010110101110010: color_data = 12'b111011101110;
20'b01010010110101110011: color_data = 12'b111011101110;
20'b01010010110101110100: color_data = 12'b111011101110;
20'b01010010110101110101: color_data = 12'b111011101110;
20'b01010010110101110110: color_data = 12'b111011101110;
20'b01010010110101110111: color_data = 12'b111011101110;
20'b01010010110101111000: color_data = 12'b111011101110;
20'b01010010110101111001: color_data = 12'b111011101110;
20'b01010010110101111011: color_data = 12'b111011101110;
20'b01010010110101111100: color_data = 12'b111011101110;
20'b01010010110101111101: color_data = 12'b111011101110;
20'b01010010110101111110: color_data = 12'b111011101110;
20'b01010010110101111111: color_data = 12'b111011101110;
20'b01010010110110000000: color_data = 12'b111011101110;
20'b01010010110110000001: color_data = 12'b111011101110;
20'b01010010110110000010: color_data = 12'b111011101110;
20'b01010010110110000011: color_data = 12'b111011101110;
20'b01010010110110000100: color_data = 12'b111011101110;
20'b01010010110110000110: color_data = 12'b111011101110;
20'b01010010110110000111: color_data = 12'b111011101110;
20'b01010010110110001000: color_data = 12'b111011101110;
20'b01010010110110001001: color_data = 12'b111011101110;
20'b01010010110110001010: color_data = 12'b111011101110;
20'b01010010110110001011: color_data = 12'b111011101110;
20'b01010010110110001100: color_data = 12'b111011101110;
20'b01010010110110001101: color_data = 12'b111011101110;
20'b01010010110110001110: color_data = 12'b111011101110;
20'b01010010110110001111: color_data = 12'b111011101110;
20'b01010010110110011100: color_data = 12'b111011101110;
20'b01010010110110011101: color_data = 12'b111011101110;
20'b01010010110110011110: color_data = 12'b111011101110;
20'b01010010110110011111: color_data = 12'b111011101110;
20'b01010010110110100000: color_data = 12'b111011101110;
20'b01010010110110100001: color_data = 12'b111011101110;
20'b01010010110110100010: color_data = 12'b111011101110;
20'b01010010110110100011: color_data = 12'b111011101110;
20'b01010010110110100100: color_data = 12'b111011101110;
20'b01010010110110100101: color_data = 12'b111011101110;
20'b01010010110110100111: color_data = 12'b111011101110;
20'b01010010110110101000: color_data = 12'b111011101110;
20'b01010010110110101001: color_data = 12'b111011101110;
20'b01010010110110101010: color_data = 12'b111011101110;
20'b01010010110110101011: color_data = 12'b111011101110;
20'b01010010110110101100: color_data = 12'b111011101110;
20'b01010010110110101101: color_data = 12'b111011101110;
20'b01010010110110101110: color_data = 12'b111011101110;
20'b01010010110110101111: color_data = 12'b111011101110;
20'b01010010110110110000: color_data = 12'b111011101110;
20'b01010010110111001000: color_data = 12'b111011101110;
20'b01010010110111001001: color_data = 12'b111011101110;
20'b01010010110111001010: color_data = 12'b111011101110;
20'b01010010110111001011: color_data = 12'b111011101110;
20'b01010010110111001100: color_data = 12'b111011101110;
20'b01010010110111001101: color_data = 12'b111011101110;
20'b01010010110111001110: color_data = 12'b111011101110;
20'b01010010110111001111: color_data = 12'b111011101110;
20'b01010010110111010000: color_data = 12'b111011101110;
20'b01010010110111010001: color_data = 12'b111011101110;
20'b01010010110111010011: color_data = 12'b111011101110;
20'b01010010110111010100: color_data = 12'b111011101110;
20'b01010010110111010101: color_data = 12'b111011101110;
20'b01010010110111010110: color_data = 12'b111011101110;
20'b01010010110111010111: color_data = 12'b111011101110;
20'b01010010110111011000: color_data = 12'b111011101110;
20'b01010010110111011001: color_data = 12'b111011101110;
20'b01010010110111011010: color_data = 12'b111011101110;
20'b01010010110111011011: color_data = 12'b111011101110;
20'b01010010110111011100: color_data = 12'b111011101110;
20'b01010011010010100001: color_data = 12'b111011101110;
20'b01010011010010100010: color_data = 12'b111011101110;
20'b01010011010010100011: color_data = 12'b111011101110;
20'b01010011010010100100: color_data = 12'b111011101110;
20'b01010011010010100101: color_data = 12'b111011101110;
20'b01010011010010100110: color_data = 12'b111011101110;
20'b01010011010010100111: color_data = 12'b111011101110;
20'b01010011010010101000: color_data = 12'b111011101110;
20'b01010011010010101001: color_data = 12'b111011101110;
20'b01010011010010101010: color_data = 12'b111011101110;
20'b01010011010010101100: color_data = 12'b111011101110;
20'b01010011010010101101: color_data = 12'b111011101110;
20'b01010011010010101110: color_data = 12'b111011101110;
20'b01010011010010101111: color_data = 12'b111011101110;
20'b01010011010010110000: color_data = 12'b111011101110;
20'b01010011010010110001: color_data = 12'b111011101110;
20'b01010011010010110010: color_data = 12'b111011101110;
20'b01010011010010110011: color_data = 12'b111011101110;
20'b01010011010010110100: color_data = 12'b111011101110;
20'b01010011010010110101: color_data = 12'b111011101110;
20'b01010011010010110111: color_data = 12'b111011101110;
20'b01010011010010111000: color_data = 12'b111011101110;
20'b01010011010010111001: color_data = 12'b111011101110;
20'b01010011010010111010: color_data = 12'b111011101110;
20'b01010011010010111011: color_data = 12'b111011101110;
20'b01010011010010111100: color_data = 12'b111011101110;
20'b01010011010010111101: color_data = 12'b111011101110;
20'b01010011010010111110: color_data = 12'b111011101110;
20'b01010011010010111111: color_data = 12'b111011101110;
20'b01010011010011000000: color_data = 12'b111011101110;
20'b01010011010011000010: color_data = 12'b111011101110;
20'b01010011010011000011: color_data = 12'b111011101110;
20'b01010011010011000100: color_data = 12'b111011101110;
20'b01010011010011000101: color_data = 12'b111011101110;
20'b01010011010011000110: color_data = 12'b111011101110;
20'b01010011010011000111: color_data = 12'b111011101110;
20'b01010011010011001000: color_data = 12'b111011101110;
20'b01010011010011001001: color_data = 12'b111011101110;
20'b01010011010011001010: color_data = 12'b111011101110;
20'b01010011010011001011: color_data = 12'b111011101110;
20'b01010011010011001101: color_data = 12'b111011101110;
20'b01010011010011001110: color_data = 12'b111011101110;
20'b01010011010011001111: color_data = 12'b111011101110;
20'b01010011010011010000: color_data = 12'b111011101110;
20'b01010011010011010001: color_data = 12'b111011101110;
20'b01010011010011010010: color_data = 12'b111011101110;
20'b01010011010011010011: color_data = 12'b111011101110;
20'b01010011010011010100: color_data = 12'b111011101110;
20'b01010011010011010101: color_data = 12'b111011101110;
20'b01010011010011010110: color_data = 12'b111011101110;
20'b01010011010100000011: color_data = 12'b111011101110;
20'b01010011010100000100: color_data = 12'b111011101110;
20'b01010011010100000101: color_data = 12'b111011101110;
20'b01010011010100000110: color_data = 12'b111011101110;
20'b01010011010100000111: color_data = 12'b111011101110;
20'b01010011010100001000: color_data = 12'b111011101110;
20'b01010011010100001001: color_data = 12'b111011101110;
20'b01010011010100001010: color_data = 12'b111011101110;
20'b01010011010100001011: color_data = 12'b111011101110;
20'b01010011010100001100: color_data = 12'b111011101110;
20'b01010011010100001110: color_data = 12'b111011101110;
20'b01010011010100001111: color_data = 12'b111011101110;
20'b01010011010100010000: color_data = 12'b111011101110;
20'b01010011010100010001: color_data = 12'b111011101110;
20'b01010011010100010010: color_data = 12'b111011101110;
20'b01010011010100010011: color_data = 12'b111011101110;
20'b01010011010100010100: color_data = 12'b111011101110;
20'b01010011010100010101: color_data = 12'b111011101110;
20'b01010011010100010110: color_data = 12'b111011101110;
20'b01010011010100010111: color_data = 12'b111011101110;
20'b01010011010100011001: color_data = 12'b111011101110;
20'b01010011010100011010: color_data = 12'b111011101110;
20'b01010011010100011011: color_data = 12'b111011101110;
20'b01010011010100011100: color_data = 12'b111011101110;
20'b01010011010100011101: color_data = 12'b111011101110;
20'b01010011010100011110: color_data = 12'b111011101110;
20'b01010011010100011111: color_data = 12'b111011101110;
20'b01010011010100100000: color_data = 12'b111011101110;
20'b01010011010100100001: color_data = 12'b111011101110;
20'b01010011010100100010: color_data = 12'b111011101110;
20'b01010011010101000100: color_data = 12'b111011101110;
20'b01010011010101000101: color_data = 12'b111011101110;
20'b01010011010101000110: color_data = 12'b111011101110;
20'b01010011010101000111: color_data = 12'b111011101110;
20'b01010011010101001000: color_data = 12'b111011101110;
20'b01010011010101001001: color_data = 12'b111011101110;
20'b01010011010101001010: color_data = 12'b111011101110;
20'b01010011010101001011: color_data = 12'b111011101110;
20'b01010011010101001100: color_data = 12'b111011101110;
20'b01010011010101001101: color_data = 12'b111011101110;
20'b01010011010101001111: color_data = 12'b111011101110;
20'b01010011010101010000: color_data = 12'b111011101110;
20'b01010011010101010001: color_data = 12'b111011101110;
20'b01010011010101010010: color_data = 12'b111011101110;
20'b01010011010101010011: color_data = 12'b111011101110;
20'b01010011010101010100: color_data = 12'b111011101110;
20'b01010011010101010101: color_data = 12'b111011101110;
20'b01010011010101010110: color_data = 12'b111011101110;
20'b01010011010101010111: color_data = 12'b111011101110;
20'b01010011010101011000: color_data = 12'b111011101110;
20'b01010011010101011010: color_data = 12'b111011101110;
20'b01010011010101011011: color_data = 12'b111011101110;
20'b01010011010101011100: color_data = 12'b111011101110;
20'b01010011010101011101: color_data = 12'b111011101110;
20'b01010011010101011110: color_data = 12'b111011101110;
20'b01010011010101011111: color_data = 12'b111011101110;
20'b01010011010101100000: color_data = 12'b111011101110;
20'b01010011010101100001: color_data = 12'b111011101110;
20'b01010011010101100010: color_data = 12'b111011101110;
20'b01010011010101100011: color_data = 12'b111011101110;
20'b01010011010101100101: color_data = 12'b111011101110;
20'b01010011010101100110: color_data = 12'b111011101110;
20'b01010011010101100111: color_data = 12'b111011101110;
20'b01010011010101101000: color_data = 12'b111011101110;
20'b01010011010101101001: color_data = 12'b111011101110;
20'b01010011010101101010: color_data = 12'b111011101110;
20'b01010011010101101011: color_data = 12'b111011101110;
20'b01010011010101101100: color_data = 12'b111011101110;
20'b01010011010101101101: color_data = 12'b111011101110;
20'b01010011010101101110: color_data = 12'b111011101110;
20'b01010011010101110000: color_data = 12'b111011101110;
20'b01010011010101110001: color_data = 12'b111011101110;
20'b01010011010101110010: color_data = 12'b111011101110;
20'b01010011010101110011: color_data = 12'b111011101110;
20'b01010011010101110100: color_data = 12'b111011101110;
20'b01010011010101110101: color_data = 12'b111011101110;
20'b01010011010101110110: color_data = 12'b111011101110;
20'b01010011010101110111: color_data = 12'b111011101110;
20'b01010011010101111000: color_data = 12'b111011101110;
20'b01010011010101111001: color_data = 12'b111011101110;
20'b01010011010101111011: color_data = 12'b111011101110;
20'b01010011010101111100: color_data = 12'b111011101110;
20'b01010011010101111101: color_data = 12'b111011101110;
20'b01010011010101111110: color_data = 12'b111011101110;
20'b01010011010101111111: color_data = 12'b111011101110;
20'b01010011010110000000: color_data = 12'b111011101110;
20'b01010011010110000001: color_data = 12'b111011101110;
20'b01010011010110000010: color_data = 12'b111011101110;
20'b01010011010110000011: color_data = 12'b111011101110;
20'b01010011010110000100: color_data = 12'b111011101110;
20'b01010011010110000110: color_data = 12'b111011101110;
20'b01010011010110000111: color_data = 12'b111011101110;
20'b01010011010110001000: color_data = 12'b111011101110;
20'b01010011010110001001: color_data = 12'b111011101110;
20'b01010011010110001010: color_data = 12'b111011101110;
20'b01010011010110001011: color_data = 12'b111011101110;
20'b01010011010110001100: color_data = 12'b111011101110;
20'b01010011010110001101: color_data = 12'b111011101110;
20'b01010011010110001110: color_data = 12'b111011101110;
20'b01010011010110001111: color_data = 12'b111011101110;
20'b01010011010110011100: color_data = 12'b111011101110;
20'b01010011010110011101: color_data = 12'b111011101110;
20'b01010011010110011110: color_data = 12'b111011101110;
20'b01010011010110011111: color_data = 12'b111011101110;
20'b01010011010110100000: color_data = 12'b111011101110;
20'b01010011010110100001: color_data = 12'b111011101110;
20'b01010011010110100010: color_data = 12'b111011101110;
20'b01010011010110100011: color_data = 12'b111011101110;
20'b01010011010110100100: color_data = 12'b111011101110;
20'b01010011010110100101: color_data = 12'b111011101110;
20'b01010011010110100111: color_data = 12'b111011101110;
20'b01010011010110101000: color_data = 12'b111011101110;
20'b01010011010110101001: color_data = 12'b111011101110;
20'b01010011010110101010: color_data = 12'b111011101110;
20'b01010011010110101011: color_data = 12'b111011101110;
20'b01010011010110101100: color_data = 12'b111011101110;
20'b01010011010110101101: color_data = 12'b111011101110;
20'b01010011010110101110: color_data = 12'b111011101110;
20'b01010011010110101111: color_data = 12'b111011101110;
20'b01010011010110110000: color_data = 12'b111011101110;
20'b01010011010111010011: color_data = 12'b111011101110;
20'b01010011010111010100: color_data = 12'b111011101110;
20'b01010011010111010101: color_data = 12'b111011101110;
20'b01010011010111010110: color_data = 12'b111011101110;
20'b01010011010111010111: color_data = 12'b111011101110;
20'b01010011010111011000: color_data = 12'b111011101110;
20'b01010011010111011001: color_data = 12'b111011101110;
20'b01010011010111011010: color_data = 12'b111011101110;
20'b01010011010111011011: color_data = 12'b111011101110;
20'b01010011010111011100: color_data = 12'b111011101110;
20'b01010011010111011110: color_data = 12'b111011101110;
20'b01010011010111011111: color_data = 12'b111011101110;
20'b01010011010111100000: color_data = 12'b111011101110;
20'b01010011010111100001: color_data = 12'b111011101110;
20'b01010011010111100010: color_data = 12'b111011101110;
20'b01010011010111100011: color_data = 12'b111011101110;
20'b01010011010111100100: color_data = 12'b111011101110;
20'b01010011010111100101: color_data = 12'b111011101110;
20'b01010011010111100110: color_data = 12'b111011101110;
20'b01010011010111100111: color_data = 12'b111011101110;
20'b01010011100010100001: color_data = 12'b111011101110;
20'b01010011100010100010: color_data = 12'b111011101110;
20'b01010011100010100011: color_data = 12'b111011101110;
20'b01010011100010100100: color_data = 12'b111011101110;
20'b01010011100010100101: color_data = 12'b111011101110;
20'b01010011100010100110: color_data = 12'b111011101110;
20'b01010011100010100111: color_data = 12'b111011101110;
20'b01010011100010101000: color_data = 12'b111011101110;
20'b01010011100010101001: color_data = 12'b111011101110;
20'b01010011100010101010: color_data = 12'b111011101110;
20'b01010011100010101100: color_data = 12'b111011101110;
20'b01010011100010101101: color_data = 12'b111011101110;
20'b01010011100010101110: color_data = 12'b111011101110;
20'b01010011100010101111: color_data = 12'b111011101110;
20'b01010011100010110000: color_data = 12'b111011101110;
20'b01010011100010110001: color_data = 12'b111011101110;
20'b01010011100010110010: color_data = 12'b111011101110;
20'b01010011100010110011: color_data = 12'b111011101110;
20'b01010011100010110100: color_data = 12'b111011101110;
20'b01010011100010110101: color_data = 12'b111011101110;
20'b01010011100010110111: color_data = 12'b111011101110;
20'b01010011100010111000: color_data = 12'b111011101110;
20'b01010011100010111001: color_data = 12'b111011101110;
20'b01010011100010111010: color_data = 12'b111011101110;
20'b01010011100010111011: color_data = 12'b111011101110;
20'b01010011100010111100: color_data = 12'b111011101110;
20'b01010011100010111101: color_data = 12'b111011101110;
20'b01010011100010111110: color_data = 12'b111011101110;
20'b01010011100010111111: color_data = 12'b111011101110;
20'b01010011100011000000: color_data = 12'b111011101110;
20'b01010011100011000010: color_data = 12'b111011101110;
20'b01010011100011000011: color_data = 12'b111011101110;
20'b01010011100011000100: color_data = 12'b111011101110;
20'b01010011100011000101: color_data = 12'b111011101110;
20'b01010011100011000110: color_data = 12'b111011101110;
20'b01010011100011000111: color_data = 12'b111011101110;
20'b01010011100011001000: color_data = 12'b111011101110;
20'b01010011100011001001: color_data = 12'b111011101110;
20'b01010011100011001010: color_data = 12'b111011101110;
20'b01010011100011001011: color_data = 12'b111011101110;
20'b01010011100011001101: color_data = 12'b111011101110;
20'b01010011100011001110: color_data = 12'b111011101110;
20'b01010011100011001111: color_data = 12'b111011101110;
20'b01010011100011010000: color_data = 12'b111011101110;
20'b01010011100011010001: color_data = 12'b111011101110;
20'b01010011100011010010: color_data = 12'b111011101110;
20'b01010011100011010011: color_data = 12'b111011101110;
20'b01010011100011010100: color_data = 12'b111011101110;
20'b01010011100011010101: color_data = 12'b111011101110;
20'b01010011100011010110: color_data = 12'b111011101110;
20'b01010011100100000011: color_data = 12'b111011101110;
20'b01010011100100000100: color_data = 12'b111011101110;
20'b01010011100100000101: color_data = 12'b111011101110;
20'b01010011100100000110: color_data = 12'b111011101110;
20'b01010011100100000111: color_data = 12'b111011101110;
20'b01010011100100001000: color_data = 12'b111011101110;
20'b01010011100100001001: color_data = 12'b111011101110;
20'b01010011100100001010: color_data = 12'b111011101110;
20'b01010011100100001011: color_data = 12'b111011101110;
20'b01010011100100001100: color_data = 12'b111011101110;
20'b01010011100100001110: color_data = 12'b111011101110;
20'b01010011100100001111: color_data = 12'b111011101110;
20'b01010011100100010000: color_data = 12'b111011101110;
20'b01010011100100010001: color_data = 12'b111011101110;
20'b01010011100100010010: color_data = 12'b111011101110;
20'b01010011100100010011: color_data = 12'b111011101110;
20'b01010011100100010100: color_data = 12'b111011101110;
20'b01010011100100010101: color_data = 12'b111011101110;
20'b01010011100100010110: color_data = 12'b111011101110;
20'b01010011100100010111: color_data = 12'b111011101110;
20'b01010011100100011001: color_data = 12'b111011101110;
20'b01010011100100011010: color_data = 12'b111011101110;
20'b01010011100100011011: color_data = 12'b111011101110;
20'b01010011100100011100: color_data = 12'b111011101110;
20'b01010011100100011101: color_data = 12'b111011101110;
20'b01010011100100011110: color_data = 12'b111011101110;
20'b01010011100100011111: color_data = 12'b111011101110;
20'b01010011100100100000: color_data = 12'b111011101110;
20'b01010011100100100001: color_data = 12'b111011101110;
20'b01010011100100100010: color_data = 12'b111011101110;
20'b01010011100101000100: color_data = 12'b111011101110;
20'b01010011100101000101: color_data = 12'b111011101110;
20'b01010011100101000110: color_data = 12'b111011101110;
20'b01010011100101000111: color_data = 12'b111011101110;
20'b01010011100101001000: color_data = 12'b111011101110;
20'b01010011100101001001: color_data = 12'b111011101110;
20'b01010011100101001010: color_data = 12'b111011101110;
20'b01010011100101001011: color_data = 12'b111011101110;
20'b01010011100101001100: color_data = 12'b111011101110;
20'b01010011100101001101: color_data = 12'b111011101110;
20'b01010011100101001111: color_data = 12'b111011101110;
20'b01010011100101010000: color_data = 12'b111011101110;
20'b01010011100101010001: color_data = 12'b111011101110;
20'b01010011100101010010: color_data = 12'b111011101110;
20'b01010011100101010011: color_data = 12'b111011101110;
20'b01010011100101010100: color_data = 12'b111011101110;
20'b01010011100101010101: color_data = 12'b111011101110;
20'b01010011100101010110: color_data = 12'b111011101110;
20'b01010011100101010111: color_data = 12'b111011101110;
20'b01010011100101011000: color_data = 12'b111011101110;
20'b01010011100101011010: color_data = 12'b111011101110;
20'b01010011100101011011: color_data = 12'b111011101110;
20'b01010011100101011100: color_data = 12'b111011101110;
20'b01010011100101011101: color_data = 12'b111011101110;
20'b01010011100101011110: color_data = 12'b111011101110;
20'b01010011100101011111: color_data = 12'b111011101110;
20'b01010011100101100000: color_data = 12'b111011101110;
20'b01010011100101100001: color_data = 12'b111011101110;
20'b01010011100101100010: color_data = 12'b111011101110;
20'b01010011100101100011: color_data = 12'b111011101110;
20'b01010011100101100101: color_data = 12'b111011101110;
20'b01010011100101100110: color_data = 12'b111011101110;
20'b01010011100101100111: color_data = 12'b111011101110;
20'b01010011100101101000: color_data = 12'b111011101110;
20'b01010011100101101001: color_data = 12'b111011101110;
20'b01010011100101101010: color_data = 12'b111011101110;
20'b01010011100101101011: color_data = 12'b111011101110;
20'b01010011100101101100: color_data = 12'b111011101110;
20'b01010011100101101101: color_data = 12'b111011101110;
20'b01010011100101101110: color_data = 12'b111011101110;
20'b01010011100101110000: color_data = 12'b111011101110;
20'b01010011100101110001: color_data = 12'b111011101110;
20'b01010011100101110010: color_data = 12'b111011101110;
20'b01010011100101110011: color_data = 12'b111011101110;
20'b01010011100101110100: color_data = 12'b111011101110;
20'b01010011100101110101: color_data = 12'b111011101110;
20'b01010011100101110110: color_data = 12'b111011101110;
20'b01010011100101110111: color_data = 12'b111011101110;
20'b01010011100101111000: color_data = 12'b111011101110;
20'b01010011100101111001: color_data = 12'b111011101110;
20'b01010011100101111011: color_data = 12'b111011101110;
20'b01010011100101111100: color_data = 12'b111011101110;
20'b01010011100101111101: color_data = 12'b111011101110;
20'b01010011100101111110: color_data = 12'b111011101110;
20'b01010011100101111111: color_data = 12'b111011101110;
20'b01010011100110000000: color_data = 12'b111011101110;
20'b01010011100110000001: color_data = 12'b111011101110;
20'b01010011100110000010: color_data = 12'b111011101110;
20'b01010011100110000011: color_data = 12'b111011101110;
20'b01010011100110000100: color_data = 12'b111011101110;
20'b01010011100110000110: color_data = 12'b111011101110;
20'b01010011100110000111: color_data = 12'b111011101110;
20'b01010011100110001000: color_data = 12'b111011101110;
20'b01010011100110001001: color_data = 12'b111011101110;
20'b01010011100110001010: color_data = 12'b111011101110;
20'b01010011100110001011: color_data = 12'b111011101110;
20'b01010011100110001100: color_data = 12'b111011101110;
20'b01010011100110001101: color_data = 12'b111011101110;
20'b01010011100110001110: color_data = 12'b111011101110;
20'b01010011100110001111: color_data = 12'b111011101110;
20'b01010011100110011100: color_data = 12'b111011101110;
20'b01010011100110011101: color_data = 12'b111011101110;
20'b01010011100110011110: color_data = 12'b111011101110;
20'b01010011100110011111: color_data = 12'b111011101110;
20'b01010011100110100000: color_data = 12'b111011101110;
20'b01010011100110100001: color_data = 12'b111011101110;
20'b01010011100110100010: color_data = 12'b111011101110;
20'b01010011100110100011: color_data = 12'b111011101110;
20'b01010011100110100100: color_data = 12'b111011101110;
20'b01010011100110100101: color_data = 12'b111011101110;
20'b01010011100110100111: color_data = 12'b111011101110;
20'b01010011100110101000: color_data = 12'b111011101110;
20'b01010011100110101001: color_data = 12'b111011101110;
20'b01010011100110101010: color_data = 12'b111011101110;
20'b01010011100110101011: color_data = 12'b111011101110;
20'b01010011100110101100: color_data = 12'b111011101110;
20'b01010011100110101101: color_data = 12'b111011101110;
20'b01010011100110101110: color_data = 12'b111011101110;
20'b01010011100110101111: color_data = 12'b111011101110;
20'b01010011100110110000: color_data = 12'b111011101110;
20'b01010011100111010011: color_data = 12'b111011101110;
20'b01010011100111010100: color_data = 12'b111011101110;
20'b01010011100111010101: color_data = 12'b111011101110;
20'b01010011100111010110: color_data = 12'b111011101110;
20'b01010011100111010111: color_data = 12'b111011101110;
20'b01010011100111011000: color_data = 12'b111011101110;
20'b01010011100111011001: color_data = 12'b111011101110;
20'b01010011100111011010: color_data = 12'b111011101110;
20'b01010011100111011011: color_data = 12'b111011101110;
20'b01010011100111011100: color_data = 12'b111011101110;
20'b01010011100111011110: color_data = 12'b111011101110;
20'b01010011100111011111: color_data = 12'b111011101110;
20'b01010011100111100000: color_data = 12'b111011101110;
20'b01010011100111100001: color_data = 12'b111011101110;
20'b01010011100111100010: color_data = 12'b111011101110;
20'b01010011100111100011: color_data = 12'b111011101110;
20'b01010011100111100100: color_data = 12'b111011101110;
20'b01010011100111100101: color_data = 12'b111011101110;
20'b01010011100111100110: color_data = 12'b111011101110;
20'b01010011100111100111: color_data = 12'b111011101110;
20'b01010011110010100001: color_data = 12'b111011101110;
20'b01010011110010100010: color_data = 12'b111011101110;
20'b01010011110010100011: color_data = 12'b111011101110;
20'b01010011110010100100: color_data = 12'b111011101110;
20'b01010011110010100101: color_data = 12'b111011101110;
20'b01010011110010100110: color_data = 12'b111011101110;
20'b01010011110010100111: color_data = 12'b111011101110;
20'b01010011110010101000: color_data = 12'b111011101110;
20'b01010011110010101001: color_data = 12'b111011101110;
20'b01010011110010101010: color_data = 12'b111011101110;
20'b01010011110010101100: color_data = 12'b111011101110;
20'b01010011110010101101: color_data = 12'b111011101110;
20'b01010011110010101110: color_data = 12'b111011101110;
20'b01010011110010101111: color_data = 12'b111011101110;
20'b01010011110010110000: color_data = 12'b111011101110;
20'b01010011110010110001: color_data = 12'b111011101110;
20'b01010011110010110010: color_data = 12'b111011101110;
20'b01010011110010110011: color_data = 12'b111011101110;
20'b01010011110010110100: color_data = 12'b111011101110;
20'b01010011110010110101: color_data = 12'b111011101110;
20'b01010011110010110111: color_data = 12'b111011101110;
20'b01010011110010111000: color_data = 12'b111011101110;
20'b01010011110010111001: color_data = 12'b111011101110;
20'b01010011110010111010: color_data = 12'b111011101110;
20'b01010011110010111011: color_data = 12'b111011101110;
20'b01010011110010111100: color_data = 12'b111011101110;
20'b01010011110010111101: color_data = 12'b111011101110;
20'b01010011110010111110: color_data = 12'b111011101110;
20'b01010011110010111111: color_data = 12'b111011101110;
20'b01010011110011000000: color_data = 12'b111011101110;
20'b01010011110011000010: color_data = 12'b111011101110;
20'b01010011110011000011: color_data = 12'b111011101110;
20'b01010011110011000100: color_data = 12'b111011101110;
20'b01010011110011000101: color_data = 12'b111011101110;
20'b01010011110011000110: color_data = 12'b111011101110;
20'b01010011110011000111: color_data = 12'b111011101110;
20'b01010011110011001000: color_data = 12'b111011101110;
20'b01010011110011001001: color_data = 12'b111011101110;
20'b01010011110011001010: color_data = 12'b111011101110;
20'b01010011110011001011: color_data = 12'b111011101110;
20'b01010011110011001101: color_data = 12'b111011101110;
20'b01010011110011001110: color_data = 12'b111011101110;
20'b01010011110011001111: color_data = 12'b111011101110;
20'b01010011110011010000: color_data = 12'b111011101110;
20'b01010011110011010001: color_data = 12'b111011101110;
20'b01010011110011010010: color_data = 12'b111011101110;
20'b01010011110011010011: color_data = 12'b111011101110;
20'b01010011110011010100: color_data = 12'b111011101110;
20'b01010011110011010101: color_data = 12'b111011101110;
20'b01010011110011010110: color_data = 12'b111011101110;
20'b01010011110100000011: color_data = 12'b111011101110;
20'b01010011110100000100: color_data = 12'b111011101110;
20'b01010011110100000101: color_data = 12'b111011101110;
20'b01010011110100000110: color_data = 12'b111011101110;
20'b01010011110100000111: color_data = 12'b111011101110;
20'b01010011110100001000: color_data = 12'b111011101110;
20'b01010011110100001001: color_data = 12'b111011101110;
20'b01010011110100001010: color_data = 12'b111011101110;
20'b01010011110100001011: color_data = 12'b111011101110;
20'b01010011110100001100: color_data = 12'b111011101110;
20'b01010011110100001110: color_data = 12'b111011101110;
20'b01010011110100001111: color_data = 12'b111011101110;
20'b01010011110100010000: color_data = 12'b111011101110;
20'b01010011110100010001: color_data = 12'b111011101110;
20'b01010011110100010010: color_data = 12'b111011101110;
20'b01010011110100010011: color_data = 12'b111011101110;
20'b01010011110100010100: color_data = 12'b111011101110;
20'b01010011110100010101: color_data = 12'b111011101110;
20'b01010011110100010110: color_data = 12'b111011101110;
20'b01010011110100010111: color_data = 12'b111011101110;
20'b01010011110100011001: color_data = 12'b111011101110;
20'b01010011110100011010: color_data = 12'b111011101110;
20'b01010011110100011011: color_data = 12'b111011101110;
20'b01010011110100011100: color_data = 12'b111011101110;
20'b01010011110100011101: color_data = 12'b111011101110;
20'b01010011110100011110: color_data = 12'b111011101110;
20'b01010011110100011111: color_data = 12'b111011101110;
20'b01010011110100100000: color_data = 12'b111011101110;
20'b01010011110100100001: color_data = 12'b111011101110;
20'b01010011110100100010: color_data = 12'b111011101110;
20'b01010011110101000100: color_data = 12'b111011101110;
20'b01010011110101000101: color_data = 12'b111011101110;
20'b01010011110101000110: color_data = 12'b111011101110;
20'b01010011110101000111: color_data = 12'b111011101110;
20'b01010011110101001000: color_data = 12'b111011101110;
20'b01010011110101001001: color_data = 12'b111011101110;
20'b01010011110101001010: color_data = 12'b111011101110;
20'b01010011110101001011: color_data = 12'b111011101110;
20'b01010011110101001100: color_data = 12'b111011101110;
20'b01010011110101001101: color_data = 12'b111011101110;
20'b01010011110101001111: color_data = 12'b111011101110;
20'b01010011110101010000: color_data = 12'b111011101110;
20'b01010011110101010001: color_data = 12'b111011101110;
20'b01010011110101010010: color_data = 12'b111011101110;
20'b01010011110101010011: color_data = 12'b111011101110;
20'b01010011110101010100: color_data = 12'b111011101110;
20'b01010011110101010101: color_data = 12'b111011101110;
20'b01010011110101010110: color_data = 12'b111011101110;
20'b01010011110101010111: color_data = 12'b111011101110;
20'b01010011110101011000: color_data = 12'b111011101110;
20'b01010011110101011010: color_data = 12'b111011101110;
20'b01010011110101011011: color_data = 12'b111011101110;
20'b01010011110101011100: color_data = 12'b111011101110;
20'b01010011110101011101: color_data = 12'b111011101110;
20'b01010011110101011110: color_data = 12'b111011101110;
20'b01010011110101011111: color_data = 12'b111011101110;
20'b01010011110101100000: color_data = 12'b111011101110;
20'b01010011110101100001: color_data = 12'b111011101110;
20'b01010011110101100010: color_data = 12'b111011101110;
20'b01010011110101100011: color_data = 12'b111011101110;
20'b01010011110101100101: color_data = 12'b111011101110;
20'b01010011110101100110: color_data = 12'b111011101110;
20'b01010011110101100111: color_data = 12'b111011101110;
20'b01010011110101101000: color_data = 12'b111011101110;
20'b01010011110101101001: color_data = 12'b111011101110;
20'b01010011110101101010: color_data = 12'b111011101110;
20'b01010011110101101011: color_data = 12'b111011101110;
20'b01010011110101101100: color_data = 12'b111011101110;
20'b01010011110101101101: color_data = 12'b111011101110;
20'b01010011110101101110: color_data = 12'b111011101110;
20'b01010011110101110000: color_data = 12'b111011101110;
20'b01010011110101110001: color_data = 12'b111011101110;
20'b01010011110101110010: color_data = 12'b111011101110;
20'b01010011110101110011: color_data = 12'b111011101110;
20'b01010011110101110100: color_data = 12'b111011101110;
20'b01010011110101110101: color_data = 12'b111011101110;
20'b01010011110101110110: color_data = 12'b111011101110;
20'b01010011110101110111: color_data = 12'b111011101110;
20'b01010011110101111000: color_data = 12'b111011101110;
20'b01010011110101111001: color_data = 12'b111011101110;
20'b01010011110101111011: color_data = 12'b111011101110;
20'b01010011110101111100: color_data = 12'b111011101110;
20'b01010011110101111101: color_data = 12'b111011101110;
20'b01010011110101111110: color_data = 12'b111011101110;
20'b01010011110101111111: color_data = 12'b111011101110;
20'b01010011110110000000: color_data = 12'b111011101110;
20'b01010011110110000001: color_data = 12'b111011101110;
20'b01010011110110000010: color_data = 12'b111011101110;
20'b01010011110110000011: color_data = 12'b111011101110;
20'b01010011110110000100: color_data = 12'b111011101110;
20'b01010011110110000110: color_data = 12'b111011101110;
20'b01010011110110000111: color_data = 12'b111011101110;
20'b01010011110110001000: color_data = 12'b111011101110;
20'b01010011110110001001: color_data = 12'b111011101110;
20'b01010011110110001010: color_data = 12'b111011101110;
20'b01010011110110001011: color_data = 12'b111011101110;
20'b01010011110110001100: color_data = 12'b111011101110;
20'b01010011110110001101: color_data = 12'b111011101110;
20'b01010011110110001110: color_data = 12'b111011101110;
20'b01010011110110001111: color_data = 12'b111011101110;
20'b01010011110110011100: color_data = 12'b111011101110;
20'b01010011110110011101: color_data = 12'b111011101110;
20'b01010011110110011110: color_data = 12'b111011101110;
20'b01010011110110011111: color_data = 12'b111011101110;
20'b01010011110110100000: color_data = 12'b111011101110;
20'b01010011110110100001: color_data = 12'b111011101110;
20'b01010011110110100010: color_data = 12'b111011101110;
20'b01010011110110100011: color_data = 12'b111011101110;
20'b01010011110110100100: color_data = 12'b111011101110;
20'b01010011110110100101: color_data = 12'b111011101110;
20'b01010011110110100111: color_data = 12'b111011101110;
20'b01010011110110101000: color_data = 12'b111011101110;
20'b01010011110110101001: color_data = 12'b111011101110;
20'b01010011110110101010: color_data = 12'b111011101110;
20'b01010011110110101011: color_data = 12'b111011101110;
20'b01010011110110101100: color_data = 12'b111011101110;
20'b01010011110110101101: color_data = 12'b111011101110;
20'b01010011110110101110: color_data = 12'b111011101110;
20'b01010011110110101111: color_data = 12'b111011101110;
20'b01010011110110110000: color_data = 12'b111011101110;
20'b01010011110111010011: color_data = 12'b111011101110;
20'b01010011110111010100: color_data = 12'b111011101110;
20'b01010011110111010101: color_data = 12'b111011101110;
20'b01010011110111010110: color_data = 12'b111011101110;
20'b01010011110111010111: color_data = 12'b111011101110;
20'b01010011110111011000: color_data = 12'b111011101110;
20'b01010011110111011001: color_data = 12'b111011101110;
20'b01010011110111011010: color_data = 12'b111011101110;
20'b01010011110111011011: color_data = 12'b111011101110;
20'b01010011110111011100: color_data = 12'b111011101110;
20'b01010011110111011110: color_data = 12'b111011101110;
20'b01010011110111011111: color_data = 12'b111011101110;
20'b01010011110111100000: color_data = 12'b111011101110;
20'b01010011110111100001: color_data = 12'b111011101110;
20'b01010011110111100010: color_data = 12'b111011101110;
20'b01010011110111100011: color_data = 12'b111011101110;
20'b01010011110111100100: color_data = 12'b111011101110;
20'b01010011110111100101: color_data = 12'b111011101110;
20'b01010011110111100110: color_data = 12'b111011101110;
20'b01010011110111100111: color_data = 12'b111011101110;
20'b01010100000010100001: color_data = 12'b111011101110;
20'b01010100000010100010: color_data = 12'b111011101110;
20'b01010100000010100011: color_data = 12'b111011101110;
20'b01010100000010100100: color_data = 12'b111011101110;
20'b01010100000010100101: color_data = 12'b111011101110;
20'b01010100000010100110: color_data = 12'b111011101110;
20'b01010100000010100111: color_data = 12'b111011101110;
20'b01010100000010101000: color_data = 12'b111011101110;
20'b01010100000010101001: color_data = 12'b111011101110;
20'b01010100000010101010: color_data = 12'b111011101110;
20'b01010100000010101100: color_data = 12'b111011101110;
20'b01010100000010101101: color_data = 12'b111011101110;
20'b01010100000010101110: color_data = 12'b111011101110;
20'b01010100000010101111: color_data = 12'b111011101110;
20'b01010100000010110000: color_data = 12'b111011101110;
20'b01010100000010110001: color_data = 12'b111011101110;
20'b01010100000010110010: color_data = 12'b111011101110;
20'b01010100000010110011: color_data = 12'b111011101110;
20'b01010100000010110100: color_data = 12'b111011101110;
20'b01010100000010110101: color_data = 12'b111011101110;
20'b01010100000010110111: color_data = 12'b111011101110;
20'b01010100000010111000: color_data = 12'b111011101110;
20'b01010100000010111001: color_data = 12'b111011101110;
20'b01010100000010111010: color_data = 12'b111011101110;
20'b01010100000010111011: color_data = 12'b111011101110;
20'b01010100000010111100: color_data = 12'b111011101110;
20'b01010100000010111101: color_data = 12'b111011101110;
20'b01010100000010111110: color_data = 12'b111011101110;
20'b01010100000010111111: color_data = 12'b111011101110;
20'b01010100000011000000: color_data = 12'b111011101110;
20'b01010100000011000010: color_data = 12'b111011101110;
20'b01010100000011000011: color_data = 12'b111011101110;
20'b01010100000011000100: color_data = 12'b111011101110;
20'b01010100000011000101: color_data = 12'b111011101110;
20'b01010100000011000110: color_data = 12'b111011101110;
20'b01010100000011000111: color_data = 12'b111011101110;
20'b01010100000011001000: color_data = 12'b111011101110;
20'b01010100000011001001: color_data = 12'b111011101110;
20'b01010100000011001010: color_data = 12'b111011101110;
20'b01010100000011001011: color_data = 12'b111011101110;
20'b01010100000011001101: color_data = 12'b111011101110;
20'b01010100000011001110: color_data = 12'b111011101110;
20'b01010100000011001111: color_data = 12'b111011101110;
20'b01010100000011010000: color_data = 12'b111011101110;
20'b01010100000011010001: color_data = 12'b111011101110;
20'b01010100000011010010: color_data = 12'b111011101110;
20'b01010100000011010011: color_data = 12'b111011101110;
20'b01010100000011010100: color_data = 12'b111011101110;
20'b01010100000011010101: color_data = 12'b111011101110;
20'b01010100000011010110: color_data = 12'b111011101110;
20'b01010100000100000011: color_data = 12'b111011101110;
20'b01010100000100000100: color_data = 12'b111011101110;
20'b01010100000100000101: color_data = 12'b111011101110;
20'b01010100000100000110: color_data = 12'b111011101110;
20'b01010100000100000111: color_data = 12'b111011101110;
20'b01010100000100001000: color_data = 12'b111011101110;
20'b01010100000100001001: color_data = 12'b111011101110;
20'b01010100000100001010: color_data = 12'b111011101110;
20'b01010100000100001011: color_data = 12'b111011101110;
20'b01010100000100001100: color_data = 12'b111011101110;
20'b01010100000100001110: color_data = 12'b111011101110;
20'b01010100000100001111: color_data = 12'b111011101110;
20'b01010100000100010000: color_data = 12'b111011101110;
20'b01010100000100010001: color_data = 12'b111011101110;
20'b01010100000100010010: color_data = 12'b111011101110;
20'b01010100000100010011: color_data = 12'b111011101110;
20'b01010100000100010100: color_data = 12'b111011101110;
20'b01010100000100010101: color_data = 12'b111011101110;
20'b01010100000100010110: color_data = 12'b111011101110;
20'b01010100000100010111: color_data = 12'b111011101110;
20'b01010100000100011001: color_data = 12'b111011101110;
20'b01010100000100011010: color_data = 12'b111011101110;
20'b01010100000100011011: color_data = 12'b111011101110;
20'b01010100000100011100: color_data = 12'b111011101110;
20'b01010100000100011101: color_data = 12'b111011101110;
20'b01010100000100011110: color_data = 12'b111011101110;
20'b01010100000100011111: color_data = 12'b111011101110;
20'b01010100000100100000: color_data = 12'b111011101110;
20'b01010100000100100001: color_data = 12'b111011101110;
20'b01010100000100100010: color_data = 12'b111011101110;
20'b01010100000101000100: color_data = 12'b111011101110;
20'b01010100000101000101: color_data = 12'b111011101110;
20'b01010100000101000110: color_data = 12'b111011101110;
20'b01010100000101000111: color_data = 12'b111011101110;
20'b01010100000101001000: color_data = 12'b111011101110;
20'b01010100000101001001: color_data = 12'b111011101110;
20'b01010100000101001010: color_data = 12'b111011101110;
20'b01010100000101001011: color_data = 12'b111011101110;
20'b01010100000101001100: color_data = 12'b111011101110;
20'b01010100000101001101: color_data = 12'b111011101110;
20'b01010100000101001111: color_data = 12'b111011101110;
20'b01010100000101010000: color_data = 12'b111011101110;
20'b01010100000101010001: color_data = 12'b111011101110;
20'b01010100000101010010: color_data = 12'b111011101110;
20'b01010100000101010011: color_data = 12'b111011101110;
20'b01010100000101010100: color_data = 12'b111011101110;
20'b01010100000101010101: color_data = 12'b111011101110;
20'b01010100000101010110: color_data = 12'b111011101110;
20'b01010100000101010111: color_data = 12'b111011101110;
20'b01010100000101011000: color_data = 12'b111011101110;
20'b01010100000101011010: color_data = 12'b111011101110;
20'b01010100000101011011: color_data = 12'b111011101110;
20'b01010100000101011100: color_data = 12'b111011101110;
20'b01010100000101011101: color_data = 12'b111011101110;
20'b01010100000101011110: color_data = 12'b111011101110;
20'b01010100000101011111: color_data = 12'b111011101110;
20'b01010100000101100000: color_data = 12'b111011101110;
20'b01010100000101100001: color_data = 12'b111011101110;
20'b01010100000101100010: color_data = 12'b111011101110;
20'b01010100000101100011: color_data = 12'b111011101110;
20'b01010100000101100101: color_data = 12'b111011101110;
20'b01010100000101100110: color_data = 12'b111011101110;
20'b01010100000101100111: color_data = 12'b111011101110;
20'b01010100000101101000: color_data = 12'b111011101110;
20'b01010100000101101001: color_data = 12'b111011101110;
20'b01010100000101101010: color_data = 12'b111011101110;
20'b01010100000101101011: color_data = 12'b111011101110;
20'b01010100000101101100: color_data = 12'b111011101110;
20'b01010100000101101101: color_data = 12'b111011101110;
20'b01010100000101101110: color_data = 12'b111011101110;
20'b01010100000101110000: color_data = 12'b111011101110;
20'b01010100000101110001: color_data = 12'b111011101110;
20'b01010100000101110010: color_data = 12'b111011101110;
20'b01010100000101110011: color_data = 12'b111011101110;
20'b01010100000101110100: color_data = 12'b111011101110;
20'b01010100000101110101: color_data = 12'b111011101110;
20'b01010100000101110110: color_data = 12'b111011101110;
20'b01010100000101110111: color_data = 12'b111011101110;
20'b01010100000101111000: color_data = 12'b111011101110;
20'b01010100000101111001: color_data = 12'b111011101110;
20'b01010100000101111011: color_data = 12'b111011101110;
20'b01010100000101111100: color_data = 12'b111011101110;
20'b01010100000101111101: color_data = 12'b111011101110;
20'b01010100000101111110: color_data = 12'b111011101110;
20'b01010100000101111111: color_data = 12'b111011101110;
20'b01010100000110000000: color_data = 12'b111011101110;
20'b01010100000110000001: color_data = 12'b111011101110;
20'b01010100000110000010: color_data = 12'b111011101110;
20'b01010100000110000011: color_data = 12'b111011101110;
20'b01010100000110000100: color_data = 12'b111011101110;
20'b01010100000110000110: color_data = 12'b111011101110;
20'b01010100000110000111: color_data = 12'b111011101110;
20'b01010100000110001000: color_data = 12'b111011101110;
20'b01010100000110001001: color_data = 12'b111011101110;
20'b01010100000110001010: color_data = 12'b111011101110;
20'b01010100000110001011: color_data = 12'b111011101110;
20'b01010100000110001100: color_data = 12'b111011101110;
20'b01010100000110001101: color_data = 12'b111011101110;
20'b01010100000110001110: color_data = 12'b111011101110;
20'b01010100000110001111: color_data = 12'b111011101110;
20'b01010100000110011100: color_data = 12'b111011101110;
20'b01010100000110011101: color_data = 12'b111011101110;
20'b01010100000110011110: color_data = 12'b111011101110;
20'b01010100000110011111: color_data = 12'b111011101110;
20'b01010100000110100000: color_data = 12'b111011101110;
20'b01010100000110100001: color_data = 12'b111011101110;
20'b01010100000110100010: color_data = 12'b111011101110;
20'b01010100000110100011: color_data = 12'b111011101110;
20'b01010100000110100100: color_data = 12'b111011101110;
20'b01010100000110100101: color_data = 12'b111011101110;
20'b01010100000110100111: color_data = 12'b111011101110;
20'b01010100000110101000: color_data = 12'b111011101110;
20'b01010100000110101001: color_data = 12'b111011101110;
20'b01010100000110101010: color_data = 12'b111011101110;
20'b01010100000110101011: color_data = 12'b111011101110;
20'b01010100000110101100: color_data = 12'b111011101110;
20'b01010100000110101101: color_data = 12'b111011101110;
20'b01010100000110101110: color_data = 12'b111011101110;
20'b01010100000110101111: color_data = 12'b111011101110;
20'b01010100000110110000: color_data = 12'b111011101110;
20'b01010100000111010011: color_data = 12'b111011101110;
20'b01010100000111010100: color_data = 12'b111011101110;
20'b01010100000111010101: color_data = 12'b111011101110;
20'b01010100000111010110: color_data = 12'b111011101110;
20'b01010100000111010111: color_data = 12'b111011101110;
20'b01010100000111011000: color_data = 12'b111011101110;
20'b01010100000111011001: color_data = 12'b111011101110;
20'b01010100000111011010: color_data = 12'b111011101110;
20'b01010100000111011011: color_data = 12'b111011101110;
20'b01010100000111011100: color_data = 12'b111011101110;
20'b01010100000111011110: color_data = 12'b111011101110;
20'b01010100000111011111: color_data = 12'b111011101110;
20'b01010100000111100000: color_data = 12'b111011101110;
20'b01010100000111100001: color_data = 12'b111011101110;
20'b01010100000111100010: color_data = 12'b111011101110;
20'b01010100000111100011: color_data = 12'b111011101110;
20'b01010100000111100100: color_data = 12'b111011101110;
20'b01010100000111100101: color_data = 12'b111011101110;
20'b01010100000111100110: color_data = 12'b111011101110;
20'b01010100000111100111: color_data = 12'b111011101110;
20'b01010100010010100001: color_data = 12'b111011101110;
20'b01010100010010100010: color_data = 12'b111011101110;
20'b01010100010010100011: color_data = 12'b111011101110;
20'b01010100010010100100: color_data = 12'b111011101110;
20'b01010100010010100101: color_data = 12'b111011101110;
20'b01010100010010100110: color_data = 12'b111011101110;
20'b01010100010010100111: color_data = 12'b111011101110;
20'b01010100010010101000: color_data = 12'b111011101110;
20'b01010100010010101001: color_data = 12'b111011101110;
20'b01010100010010101010: color_data = 12'b111011101110;
20'b01010100010010101100: color_data = 12'b111011101110;
20'b01010100010010101101: color_data = 12'b111011101110;
20'b01010100010010101110: color_data = 12'b111011101110;
20'b01010100010010101111: color_data = 12'b111011101110;
20'b01010100010010110000: color_data = 12'b111011101110;
20'b01010100010010110001: color_data = 12'b111011101110;
20'b01010100010010110010: color_data = 12'b111011101110;
20'b01010100010010110011: color_data = 12'b111011101110;
20'b01010100010010110100: color_data = 12'b111011101110;
20'b01010100010010110101: color_data = 12'b111011101110;
20'b01010100010010110111: color_data = 12'b111011101110;
20'b01010100010010111000: color_data = 12'b111011101110;
20'b01010100010010111001: color_data = 12'b111011101110;
20'b01010100010010111010: color_data = 12'b111011101110;
20'b01010100010010111011: color_data = 12'b111011101110;
20'b01010100010010111100: color_data = 12'b111011101110;
20'b01010100010010111101: color_data = 12'b111011101110;
20'b01010100010010111110: color_data = 12'b111011101110;
20'b01010100010010111111: color_data = 12'b111011101110;
20'b01010100010011000000: color_data = 12'b111011101110;
20'b01010100010011000010: color_data = 12'b111011101110;
20'b01010100010011000011: color_data = 12'b111011101110;
20'b01010100010011000100: color_data = 12'b111011101110;
20'b01010100010011000101: color_data = 12'b111011101110;
20'b01010100010011000110: color_data = 12'b111011101110;
20'b01010100010011000111: color_data = 12'b111011101110;
20'b01010100010011001000: color_data = 12'b111011101110;
20'b01010100010011001001: color_data = 12'b111011101110;
20'b01010100010011001010: color_data = 12'b111011101110;
20'b01010100010011001011: color_data = 12'b111011101110;
20'b01010100010011001101: color_data = 12'b111011101110;
20'b01010100010011001110: color_data = 12'b111011101110;
20'b01010100010011001111: color_data = 12'b111011101110;
20'b01010100010011010000: color_data = 12'b111011101110;
20'b01010100010011010001: color_data = 12'b111011101110;
20'b01010100010011010010: color_data = 12'b111011101110;
20'b01010100010011010011: color_data = 12'b111011101110;
20'b01010100010011010100: color_data = 12'b111011101110;
20'b01010100010011010101: color_data = 12'b111011101110;
20'b01010100010011010110: color_data = 12'b111011101110;
20'b01010100010100000011: color_data = 12'b111011101110;
20'b01010100010100000100: color_data = 12'b111011101110;
20'b01010100010100000101: color_data = 12'b111011101110;
20'b01010100010100000110: color_data = 12'b111011101110;
20'b01010100010100000111: color_data = 12'b111011101110;
20'b01010100010100001000: color_data = 12'b111011101110;
20'b01010100010100001001: color_data = 12'b111011101110;
20'b01010100010100001010: color_data = 12'b111011101110;
20'b01010100010100001011: color_data = 12'b111011101110;
20'b01010100010100001100: color_data = 12'b111011101110;
20'b01010100010100001110: color_data = 12'b111011101110;
20'b01010100010100001111: color_data = 12'b111011101110;
20'b01010100010100010000: color_data = 12'b111011101110;
20'b01010100010100010001: color_data = 12'b111011101110;
20'b01010100010100010010: color_data = 12'b111011101110;
20'b01010100010100010011: color_data = 12'b111011101110;
20'b01010100010100010100: color_data = 12'b111011101110;
20'b01010100010100010101: color_data = 12'b111011101110;
20'b01010100010100010110: color_data = 12'b111011101110;
20'b01010100010100010111: color_data = 12'b111011101110;
20'b01010100010100011001: color_data = 12'b111011101110;
20'b01010100010100011010: color_data = 12'b111011101110;
20'b01010100010100011011: color_data = 12'b111011101110;
20'b01010100010100011100: color_data = 12'b111011101110;
20'b01010100010100011101: color_data = 12'b111011101110;
20'b01010100010100011110: color_data = 12'b111011101110;
20'b01010100010100011111: color_data = 12'b111011101110;
20'b01010100010100100000: color_data = 12'b111011101110;
20'b01010100010100100001: color_data = 12'b111011101110;
20'b01010100010100100010: color_data = 12'b111011101110;
20'b01010100010101000100: color_data = 12'b111011101110;
20'b01010100010101000101: color_data = 12'b111011101110;
20'b01010100010101000110: color_data = 12'b111011101110;
20'b01010100010101000111: color_data = 12'b111011101110;
20'b01010100010101001000: color_data = 12'b111011101110;
20'b01010100010101001001: color_data = 12'b111011101110;
20'b01010100010101001010: color_data = 12'b111011101110;
20'b01010100010101001011: color_data = 12'b111011101110;
20'b01010100010101001100: color_data = 12'b111011101110;
20'b01010100010101001101: color_data = 12'b111011101110;
20'b01010100010101001111: color_data = 12'b111011101110;
20'b01010100010101010000: color_data = 12'b111011101110;
20'b01010100010101010001: color_data = 12'b111011101110;
20'b01010100010101010010: color_data = 12'b111011101110;
20'b01010100010101010011: color_data = 12'b111011101110;
20'b01010100010101010100: color_data = 12'b111011101110;
20'b01010100010101010101: color_data = 12'b111011101110;
20'b01010100010101010110: color_data = 12'b111011101110;
20'b01010100010101010111: color_data = 12'b111011101110;
20'b01010100010101011000: color_data = 12'b111011101110;
20'b01010100010101011010: color_data = 12'b111011101110;
20'b01010100010101011011: color_data = 12'b111011101110;
20'b01010100010101011100: color_data = 12'b111011101110;
20'b01010100010101011101: color_data = 12'b111011101110;
20'b01010100010101011110: color_data = 12'b111011101110;
20'b01010100010101011111: color_data = 12'b111011101110;
20'b01010100010101100000: color_data = 12'b111011101110;
20'b01010100010101100001: color_data = 12'b111011101110;
20'b01010100010101100010: color_data = 12'b111011101110;
20'b01010100010101100011: color_data = 12'b111011101110;
20'b01010100010101100101: color_data = 12'b111011101110;
20'b01010100010101100110: color_data = 12'b111011101110;
20'b01010100010101100111: color_data = 12'b111011101110;
20'b01010100010101101000: color_data = 12'b111011101110;
20'b01010100010101101001: color_data = 12'b111011101110;
20'b01010100010101101010: color_data = 12'b111011101110;
20'b01010100010101101011: color_data = 12'b111011101110;
20'b01010100010101101100: color_data = 12'b111011101110;
20'b01010100010101101101: color_data = 12'b111011101110;
20'b01010100010101101110: color_data = 12'b111011101110;
20'b01010100010101110000: color_data = 12'b111011101110;
20'b01010100010101110001: color_data = 12'b111011101110;
20'b01010100010101110010: color_data = 12'b111011101110;
20'b01010100010101110011: color_data = 12'b111011101110;
20'b01010100010101110100: color_data = 12'b111011101110;
20'b01010100010101110101: color_data = 12'b111011101110;
20'b01010100010101110110: color_data = 12'b111011101110;
20'b01010100010101110111: color_data = 12'b111011101110;
20'b01010100010101111000: color_data = 12'b111011101110;
20'b01010100010101111001: color_data = 12'b111011101110;
20'b01010100010101111011: color_data = 12'b111011101110;
20'b01010100010101111100: color_data = 12'b111011101110;
20'b01010100010101111101: color_data = 12'b111011101110;
20'b01010100010101111110: color_data = 12'b111011101110;
20'b01010100010101111111: color_data = 12'b111011101110;
20'b01010100010110000000: color_data = 12'b111011101110;
20'b01010100010110000001: color_data = 12'b111011101110;
20'b01010100010110000010: color_data = 12'b111011101110;
20'b01010100010110000011: color_data = 12'b111011101110;
20'b01010100010110000100: color_data = 12'b111011101110;
20'b01010100010110000110: color_data = 12'b111011101110;
20'b01010100010110000111: color_data = 12'b111011101110;
20'b01010100010110001000: color_data = 12'b111011101110;
20'b01010100010110001001: color_data = 12'b111011101110;
20'b01010100010110001010: color_data = 12'b111011101110;
20'b01010100010110001011: color_data = 12'b111011101110;
20'b01010100010110001100: color_data = 12'b111011101110;
20'b01010100010110001101: color_data = 12'b111011101110;
20'b01010100010110001110: color_data = 12'b111011101110;
20'b01010100010110001111: color_data = 12'b111011101110;
20'b01010100010110011100: color_data = 12'b111011101110;
20'b01010100010110011101: color_data = 12'b111011101110;
20'b01010100010110011110: color_data = 12'b111011101110;
20'b01010100010110011111: color_data = 12'b111011101110;
20'b01010100010110100000: color_data = 12'b111011101110;
20'b01010100010110100001: color_data = 12'b111011101110;
20'b01010100010110100010: color_data = 12'b111011101110;
20'b01010100010110100011: color_data = 12'b111011101110;
20'b01010100010110100100: color_data = 12'b111011101110;
20'b01010100010110100101: color_data = 12'b111011101110;
20'b01010100010110100111: color_data = 12'b111011101110;
20'b01010100010110101000: color_data = 12'b111011101110;
20'b01010100010110101001: color_data = 12'b111011101110;
20'b01010100010110101010: color_data = 12'b111011101110;
20'b01010100010110101011: color_data = 12'b111011101110;
20'b01010100010110101100: color_data = 12'b111011101110;
20'b01010100010110101101: color_data = 12'b111011101110;
20'b01010100010110101110: color_data = 12'b111011101110;
20'b01010100010110101111: color_data = 12'b111011101110;
20'b01010100010110110000: color_data = 12'b111011101110;
20'b01010100010111010011: color_data = 12'b111011101110;
20'b01010100010111010100: color_data = 12'b111011101110;
20'b01010100010111010101: color_data = 12'b111011101110;
20'b01010100010111010110: color_data = 12'b111011101110;
20'b01010100010111010111: color_data = 12'b111011101110;
20'b01010100010111011000: color_data = 12'b111011101110;
20'b01010100010111011001: color_data = 12'b111011101110;
20'b01010100010111011010: color_data = 12'b111011101110;
20'b01010100010111011011: color_data = 12'b111011101110;
20'b01010100010111011100: color_data = 12'b111011101110;
20'b01010100010111011110: color_data = 12'b111011101110;
20'b01010100010111011111: color_data = 12'b111011101110;
20'b01010100010111100000: color_data = 12'b111011101110;
20'b01010100010111100001: color_data = 12'b111011101110;
20'b01010100010111100010: color_data = 12'b111011101110;
20'b01010100010111100011: color_data = 12'b111011101110;
20'b01010100010111100100: color_data = 12'b111011101110;
20'b01010100010111100101: color_data = 12'b111011101110;
20'b01010100010111100110: color_data = 12'b111011101110;
20'b01010100010111100111: color_data = 12'b111011101110;
20'b01010100100010100001: color_data = 12'b111011101110;
20'b01010100100010100010: color_data = 12'b111011101110;
20'b01010100100010100011: color_data = 12'b111011101110;
20'b01010100100010100100: color_data = 12'b111011101110;
20'b01010100100010100101: color_data = 12'b111011101110;
20'b01010100100010100110: color_data = 12'b111011101110;
20'b01010100100010100111: color_data = 12'b111011101110;
20'b01010100100010101000: color_data = 12'b111011101110;
20'b01010100100010101001: color_data = 12'b111011101110;
20'b01010100100010101010: color_data = 12'b111011101110;
20'b01010100100010101100: color_data = 12'b111011101110;
20'b01010100100010101101: color_data = 12'b111011101110;
20'b01010100100010101110: color_data = 12'b111011101110;
20'b01010100100010101111: color_data = 12'b111011101110;
20'b01010100100010110000: color_data = 12'b111011101110;
20'b01010100100010110001: color_data = 12'b111011101110;
20'b01010100100010110010: color_data = 12'b111011101110;
20'b01010100100010110011: color_data = 12'b111011101110;
20'b01010100100010110100: color_data = 12'b111011101110;
20'b01010100100010110101: color_data = 12'b111011101110;
20'b01010100100010110111: color_data = 12'b111011101110;
20'b01010100100010111000: color_data = 12'b111011101110;
20'b01010100100010111001: color_data = 12'b111011101110;
20'b01010100100010111010: color_data = 12'b111011101110;
20'b01010100100010111011: color_data = 12'b111011101110;
20'b01010100100010111100: color_data = 12'b111011101110;
20'b01010100100010111101: color_data = 12'b111011101110;
20'b01010100100010111110: color_data = 12'b111011101110;
20'b01010100100010111111: color_data = 12'b111011101110;
20'b01010100100011000000: color_data = 12'b111011101110;
20'b01010100100011000010: color_data = 12'b111011101110;
20'b01010100100011000011: color_data = 12'b111011101110;
20'b01010100100011000100: color_data = 12'b111011101110;
20'b01010100100011000101: color_data = 12'b111011101110;
20'b01010100100011000110: color_data = 12'b111011101110;
20'b01010100100011000111: color_data = 12'b111011101110;
20'b01010100100011001000: color_data = 12'b111011101110;
20'b01010100100011001001: color_data = 12'b111011101110;
20'b01010100100011001010: color_data = 12'b111011101110;
20'b01010100100011001011: color_data = 12'b111011101110;
20'b01010100100011001101: color_data = 12'b111011101110;
20'b01010100100011001110: color_data = 12'b111011101110;
20'b01010100100011001111: color_data = 12'b111011101110;
20'b01010100100011010000: color_data = 12'b111011101110;
20'b01010100100011010001: color_data = 12'b111011101110;
20'b01010100100011010010: color_data = 12'b111011101110;
20'b01010100100011010011: color_data = 12'b111011101110;
20'b01010100100011010100: color_data = 12'b111011101110;
20'b01010100100011010101: color_data = 12'b111011101110;
20'b01010100100011010110: color_data = 12'b111011101110;
20'b01010100100100000011: color_data = 12'b111011101110;
20'b01010100100100000100: color_data = 12'b111011101110;
20'b01010100100100000101: color_data = 12'b111011101110;
20'b01010100100100000110: color_data = 12'b111011101110;
20'b01010100100100000111: color_data = 12'b111011101110;
20'b01010100100100001000: color_data = 12'b111011101110;
20'b01010100100100001001: color_data = 12'b111011101110;
20'b01010100100100001010: color_data = 12'b111011101110;
20'b01010100100100001011: color_data = 12'b111011101110;
20'b01010100100100001100: color_data = 12'b111011101110;
20'b01010100100100001110: color_data = 12'b111011101110;
20'b01010100100100001111: color_data = 12'b111011101110;
20'b01010100100100010000: color_data = 12'b111011101110;
20'b01010100100100010001: color_data = 12'b111011101110;
20'b01010100100100010010: color_data = 12'b111011101110;
20'b01010100100100010011: color_data = 12'b111011101110;
20'b01010100100100010100: color_data = 12'b111011101110;
20'b01010100100100010101: color_data = 12'b111011101110;
20'b01010100100100010110: color_data = 12'b111011101110;
20'b01010100100100010111: color_data = 12'b111011101110;
20'b01010100100100011001: color_data = 12'b111011101110;
20'b01010100100100011010: color_data = 12'b111011101110;
20'b01010100100100011011: color_data = 12'b111011101110;
20'b01010100100100011100: color_data = 12'b111011101110;
20'b01010100100100011101: color_data = 12'b111011101110;
20'b01010100100100011110: color_data = 12'b111011101110;
20'b01010100100100011111: color_data = 12'b111011101110;
20'b01010100100100100000: color_data = 12'b111011101110;
20'b01010100100100100001: color_data = 12'b111011101110;
20'b01010100100100100010: color_data = 12'b111011101110;
20'b01010100100101000100: color_data = 12'b111011101110;
20'b01010100100101000101: color_data = 12'b111011101110;
20'b01010100100101000110: color_data = 12'b111011101110;
20'b01010100100101000111: color_data = 12'b111011101110;
20'b01010100100101001000: color_data = 12'b111011101110;
20'b01010100100101001001: color_data = 12'b111011101110;
20'b01010100100101001010: color_data = 12'b111011101110;
20'b01010100100101001011: color_data = 12'b111011101110;
20'b01010100100101001100: color_data = 12'b111011101110;
20'b01010100100101001101: color_data = 12'b111011101110;
20'b01010100100101001111: color_data = 12'b111011101110;
20'b01010100100101010000: color_data = 12'b111011101110;
20'b01010100100101010001: color_data = 12'b111011101110;
20'b01010100100101010010: color_data = 12'b111011101110;
20'b01010100100101010011: color_data = 12'b111011101110;
20'b01010100100101010100: color_data = 12'b111011101110;
20'b01010100100101010101: color_data = 12'b111011101110;
20'b01010100100101010110: color_data = 12'b111011101110;
20'b01010100100101010111: color_data = 12'b111011101110;
20'b01010100100101011000: color_data = 12'b111011101110;
20'b01010100100101011010: color_data = 12'b111011101110;
20'b01010100100101011011: color_data = 12'b111011101110;
20'b01010100100101011100: color_data = 12'b111011101110;
20'b01010100100101011101: color_data = 12'b111011101110;
20'b01010100100101011110: color_data = 12'b111011101110;
20'b01010100100101011111: color_data = 12'b111011101110;
20'b01010100100101100000: color_data = 12'b111011101110;
20'b01010100100101100001: color_data = 12'b111011101110;
20'b01010100100101100010: color_data = 12'b111011101110;
20'b01010100100101100011: color_data = 12'b111011101110;
20'b01010100100101100101: color_data = 12'b111011101110;
20'b01010100100101100110: color_data = 12'b111011101110;
20'b01010100100101100111: color_data = 12'b111011101110;
20'b01010100100101101000: color_data = 12'b111011101110;
20'b01010100100101101001: color_data = 12'b111011101110;
20'b01010100100101101010: color_data = 12'b111011101110;
20'b01010100100101101011: color_data = 12'b111011101110;
20'b01010100100101101100: color_data = 12'b111011101110;
20'b01010100100101101101: color_data = 12'b111011101110;
20'b01010100100101101110: color_data = 12'b111011101110;
20'b01010100100101110000: color_data = 12'b111011101110;
20'b01010100100101110001: color_data = 12'b111011101110;
20'b01010100100101110010: color_data = 12'b111011101110;
20'b01010100100101110011: color_data = 12'b111011101110;
20'b01010100100101110100: color_data = 12'b111011101110;
20'b01010100100101110101: color_data = 12'b111011101110;
20'b01010100100101110110: color_data = 12'b111011101110;
20'b01010100100101110111: color_data = 12'b111011101110;
20'b01010100100101111000: color_data = 12'b111011101110;
20'b01010100100101111001: color_data = 12'b111011101110;
20'b01010100100101111011: color_data = 12'b111011101110;
20'b01010100100101111100: color_data = 12'b111011101110;
20'b01010100100101111101: color_data = 12'b111011101110;
20'b01010100100101111110: color_data = 12'b111011101110;
20'b01010100100101111111: color_data = 12'b111011101110;
20'b01010100100110000000: color_data = 12'b111011101110;
20'b01010100100110000001: color_data = 12'b111011101110;
20'b01010100100110000010: color_data = 12'b111011101110;
20'b01010100100110000011: color_data = 12'b111011101110;
20'b01010100100110000100: color_data = 12'b111011101110;
20'b01010100100110000110: color_data = 12'b111011101110;
20'b01010100100110000111: color_data = 12'b111011101110;
20'b01010100100110001000: color_data = 12'b111011101110;
20'b01010100100110001001: color_data = 12'b111011101110;
20'b01010100100110001010: color_data = 12'b111011101110;
20'b01010100100110001011: color_data = 12'b111011101110;
20'b01010100100110001100: color_data = 12'b111011101110;
20'b01010100100110001101: color_data = 12'b111011101110;
20'b01010100100110001110: color_data = 12'b111011101110;
20'b01010100100110001111: color_data = 12'b111011101110;
20'b01010100100110011100: color_data = 12'b111011101110;
20'b01010100100110011101: color_data = 12'b111011101110;
20'b01010100100110011110: color_data = 12'b111011101110;
20'b01010100100110011111: color_data = 12'b111011101110;
20'b01010100100110100000: color_data = 12'b111011101110;
20'b01010100100110100001: color_data = 12'b111011101110;
20'b01010100100110100010: color_data = 12'b111011101110;
20'b01010100100110100011: color_data = 12'b111011101110;
20'b01010100100110100100: color_data = 12'b111011101110;
20'b01010100100110100101: color_data = 12'b111011101110;
20'b01010100100110100111: color_data = 12'b111011101110;
20'b01010100100110101000: color_data = 12'b111011101110;
20'b01010100100110101001: color_data = 12'b111011101110;
20'b01010100100110101010: color_data = 12'b111011101110;
20'b01010100100110101011: color_data = 12'b111011101110;
20'b01010100100110101100: color_data = 12'b111011101110;
20'b01010100100110101101: color_data = 12'b111011101110;
20'b01010100100110101110: color_data = 12'b111011101110;
20'b01010100100110101111: color_data = 12'b111011101110;
20'b01010100100110110000: color_data = 12'b111011101110;
20'b01010100100111010011: color_data = 12'b111011101110;
20'b01010100100111010100: color_data = 12'b111011101110;
20'b01010100100111010101: color_data = 12'b111011101110;
20'b01010100100111010110: color_data = 12'b111011101110;
20'b01010100100111010111: color_data = 12'b111011101110;
20'b01010100100111011000: color_data = 12'b111011101110;
20'b01010100100111011001: color_data = 12'b111011101110;
20'b01010100100111011010: color_data = 12'b111011101110;
20'b01010100100111011011: color_data = 12'b111011101110;
20'b01010100100111011100: color_data = 12'b111011101110;
20'b01010100100111011110: color_data = 12'b111011101110;
20'b01010100100111011111: color_data = 12'b111011101110;
20'b01010100100111100000: color_data = 12'b111011101110;
20'b01010100100111100001: color_data = 12'b111011101110;
20'b01010100100111100010: color_data = 12'b111011101110;
20'b01010100100111100011: color_data = 12'b111011101110;
20'b01010100100111100100: color_data = 12'b111011101110;
20'b01010100100111100101: color_data = 12'b111011101110;
20'b01010100100111100110: color_data = 12'b111011101110;
20'b01010100100111100111: color_data = 12'b111011101110;
20'b01010100110010100001: color_data = 12'b111011101110;
20'b01010100110010100010: color_data = 12'b111011101110;
20'b01010100110010100011: color_data = 12'b111011101110;
20'b01010100110010100100: color_data = 12'b111011101110;
20'b01010100110010100101: color_data = 12'b111011101110;
20'b01010100110010100110: color_data = 12'b111011101110;
20'b01010100110010100111: color_data = 12'b111011101110;
20'b01010100110010101000: color_data = 12'b111011101110;
20'b01010100110010101001: color_data = 12'b111011101110;
20'b01010100110010101010: color_data = 12'b111011101110;
20'b01010100110010101100: color_data = 12'b111011101110;
20'b01010100110010101101: color_data = 12'b111011101110;
20'b01010100110010101110: color_data = 12'b111011101110;
20'b01010100110010101111: color_data = 12'b111011101110;
20'b01010100110010110000: color_data = 12'b111011101110;
20'b01010100110010110001: color_data = 12'b111011101110;
20'b01010100110010110010: color_data = 12'b111011101110;
20'b01010100110010110011: color_data = 12'b111011101110;
20'b01010100110010110100: color_data = 12'b111011101110;
20'b01010100110010110101: color_data = 12'b111011101110;
20'b01010100110010110111: color_data = 12'b111011101110;
20'b01010100110010111000: color_data = 12'b111011101110;
20'b01010100110010111001: color_data = 12'b111011101110;
20'b01010100110010111010: color_data = 12'b111011101110;
20'b01010100110010111011: color_data = 12'b111011101110;
20'b01010100110010111100: color_data = 12'b111011101110;
20'b01010100110010111101: color_data = 12'b111011101110;
20'b01010100110010111110: color_data = 12'b111011101110;
20'b01010100110010111111: color_data = 12'b111011101110;
20'b01010100110011000000: color_data = 12'b111011101110;
20'b01010100110011000010: color_data = 12'b111011101110;
20'b01010100110011000011: color_data = 12'b111011101110;
20'b01010100110011000100: color_data = 12'b111011101110;
20'b01010100110011000101: color_data = 12'b111011101110;
20'b01010100110011000110: color_data = 12'b111011101110;
20'b01010100110011000111: color_data = 12'b111011101110;
20'b01010100110011001000: color_data = 12'b111011101110;
20'b01010100110011001001: color_data = 12'b111011101110;
20'b01010100110011001010: color_data = 12'b111011101110;
20'b01010100110011001011: color_data = 12'b111011101110;
20'b01010100110011001101: color_data = 12'b111011101110;
20'b01010100110011001110: color_data = 12'b111011101110;
20'b01010100110011001111: color_data = 12'b111011101110;
20'b01010100110011010000: color_data = 12'b111011101110;
20'b01010100110011010001: color_data = 12'b111011101110;
20'b01010100110011010010: color_data = 12'b111011101110;
20'b01010100110011010011: color_data = 12'b111011101110;
20'b01010100110011010100: color_data = 12'b111011101110;
20'b01010100110011010101: color_data = 12'b111011101110;
20'b01010100110011010110: color_data = 12'b111011101110;
20'b01010100110100000011: color_data = 12'b111011101110;
20'b01010100110100000100: color_data = 12'b111011101110;
20'b01010100110100000101: color_data = 12'b111011101110;
20'b01010100110100000110: color_data = 12'b111011101110;
20'b01010100110100000111: color_data = 12'b111011101110;
20'b01010100110100001000: color_data = 12'b111011101110;
20'b01010100110100001001: color_data = 12'b111011101110;
20'b01010100110100001010: color_data = 12'b111011101110;
20'b01010100110100001011: color_data = 12'b111011101110;
20'b01010100110100001100: color_data = 12'b111011101110;
20'b01010100110100001110: color_data = 12'b111011101110;
20'b01010100110100001111: color_data = 12'b111011101110;
20'b01010100110100010000: color_data = 12'b111011101110;
20'b01010100110100010001: color_data = 12'b111011101110;
20'b01010100110100010010: color_data = 12'b111011101110;
20'b01010100110100010011: color_data = 12'b111011101110;
20'b01010100110100010100: color_data = 12'b111011101110;
20'b01010100110100010101: color_data = 12'b111011101110;
20'b01010100110100010110: color_data = 12'b111011101110;
20'b01010100110100010111: color_data = 12'b111011101110;
20'b01010100110100011001: color_data = 12'b111011101110;
20'b01010100110100011010: color_data = 12'b111011101110;
20'b01010100110100011011: color_data = 12'b111011101110;
20'b01010100110100011100: color_data = 12'b111011101110;
20'b01010100110100011101: color_data = 12'b111011101110;
20'b01010100110100011110: color_data = 12'b111011101110;
20'b01010100110100011111: color_data = 12'b111011101110;
20'b01010100110100100000: color_data = 12'b111011101110;
20'b01010100110100100001: color_data = 12'b111011101110;
20'b01010100110100100010: color_data = 12'b111011101110;
20'b01010100110101000100: color_data = 12'b111011101110;
20'b01010100110101000101: color_data = 12'b111011101110;
20'b01010100110101000110: color_data = 12'b111011101110;
20'b01010100110101000111: color_data = 12'b111011101110;
20'b01010100110101001000: color_data = 12'b111011101110;
20'b01010100110101001001: color_data = 12'b111011101110;
20'b01010100110101001010: color_data = 12'b111011101110;
20'b01010100110101001011: color_data = 12'b111011101110;
20'b01010100110101001100: color_data = 12'b111011101110;
20'b01010100110101001101: color_data = 12'b111011101110;
20'b01010100110101001111: color_data = 12'b111011101110;
20'b01010100110101010000: color_data = 12'b111011101110;
20'b01010100110101010001: color_data = 12'b111011101110;
20'b01010100110101010010: color_data = 12'b111011101110;
20'b01010100110101010011: color_data = 12'b111011101110;
20'b01010100110101010100: color_data = 12'b111011101110;
20'b01010100110101010101: color_data = 12'b111011101110;
20'b01010100110101010110: color_data = 12'b111011101110;
20'b01010100110101010111: color_data = 12'b111011101110;
20'b01010100110101011000: color_data = 12'b111011101110;
20'b01010100110101011010: color_data = 12'b111011101110;
20'b01010100110101011011: color_data = 12'b111011101110;
20'b01010100110101011100: color_data = 12'b111011101110;
20'b01010100110101011101: color_data = 12'b111011101110;
20'b01010100110101011110: color_data = 12'b111011101110;
20'b01010100110101011111: color_data = 12'b111011101110;
20'b01010100110101100000: color_data = 12'b111011101110;
20'b01010100110101100001: color_data = 12'b111011101110;
20'b01010100110101100010: color_data = 12'b111011101110;
20'b01010100110101100011: color_data = 12'b111011101110;
20'b01010100110101100101: color_data = 12'b111011101110;
20'b01010100110101100110: color_data = 12'b111011101110;
20'b01010100110101100111: color_data = 12'b111011101110;
20'b01010100110101101000: color_data = 12'b111011101110;
20'b01010100110101101001: color_data = 12'b111011101110;
20'b01010100110101101010: color_data = 12'b111011101110;
20'b01010100110101101011: color_data = 12'b111011101110;
20'b01010100110101101100: color_data = 12'b111011101110;
20'b01010100110101101101: color_data = 12'b111011101110;
20'b01010100110101101110: color_data = 12'b111011101110;
20'b01010100110101110000: color_data = 12'b111011101110;
20'b01010100110101110001: color_data = 12'b111011101110;
20'b01010100110101110010: color_data = 12'b111011101110;
20'b01010100110101110011: color_data = 12'b111011101110;
20'b01010100110101110100: color_data = 12'b111011101110;
20'b01010100110101110101: color_data = 12'b111011101110;
20'b01010100110101110110: color_data = 12'b111011101110;
20'b01010100110101110111: color_data = 12'b111011101110;
20'b01010100110101111000: color_data = 12'b111011101110;
20'b01010100110101111001: color_data = 12'b111011101110;
20'b01010100110101111011: color_data = 12'b111011101110;
20'b01010100110101111100: color_data = 12'b111011101110;
20'b01010100110101111101: color_data = 12'b111011101110;
20'b01010100110101111110: color_data = 12'b111011101110;
20'b01010100110101111111: color_data = 12'b111011101110;
20'b01010100110110000000: color_data = 12'b111011101110;
20'b01010100110110000001: color_data = 12'b111011101110;
20'b01010100110110000010: color_data = 12'b111011101110;
20'b01010100110110000011: color_data = 12'b111011101110;
20'b01010100110110000100: color_data = 12'b111011101110;
20'b01010100110110000110: color_data = 12'b111011101110;
20'b01010100110110000111: color_data = 12'b111011101110;
20'b01010100110110001000: color_data = 12'b111011101110;
20'b01010100110110001001: color_data = 12'b111011101110;
20'b01010100110110001010: color_data = 12'b111011101110;
20'b01010100110110001011: color_data = 12'b111011101110;
20'b01010100110110001100: color_data = 12'b111011101110;
20'b01010100110110001101: color_data = 12'b111011101110;
20'b01010100110110001110: color_data = 12'b111011101110;
20'b01010100110110001111: color_data = 12'b111011101110;
20'b01010100110110011100: color_data = 12'b111011101110;
20'b01010100110110011101: color_data = 12'b111011101110;
20'b01010100110110011110: color_data = 12'b111011101110;
20'b01010100110110011111: color_data = 12'b111011101110;
20'b01010100110110100000: color_data = 12'b111011101110;
20'b01010100110110100001: color_data = 12'b111011101110;
20'b01010100110110100010: color_data = 12'b111011101110;
20'b01010100110110100011: color_data = 12'b111011101110;
20'b01010100110110100100: color_data = 12'b111011101110;
20'b01010100110110100101: color_data = 12'b111011101110;
20'b01010100110110100111: color_data = 12'b111011101110;
20'b01010100110110101000: color_data = 12'b111011101110;
20'b01010100110110101001: color_data = 12'b111011101110;
20'b01010100110110101010: color_data = 12'b111011101110;
20'b01010100110110101011: color_data = 12'b111011101110;
20'b01010100110110101100: color_data = 12'b111011101110;
20'b01010100110110101101: color_data = 12'b111011101110;
20'b01010100110110101110: color_data = 12'b111011101110;
20'b01010100110110101111: color_data = 12'b111011101110;
20'b01010100110110110000: color_data = 12'b111011101110;
20'b01010100110111010011: color_data = 12'b111011101110;
20'b01010100110111010100: color_data = 12'b111011101110;
20'b01010100110111010101: color_data = 12'b111011101110;
20'b01010100110111010110: color_data = 12'b111011101110;
20'b01010100110111010111: color_data = 12'b111011101110;
20'b01010100110111011000: color_data = 12'b111011101110;
20'b01010100110111011001: color_data = 12'b111011101110;
20'b01010100110111011010: color_data = 12'b111011101110;
20'b01010100110111011011: color_data = 12'b111011101110;
20'b01010100110111011100: color_data = 12'b111011101110;
20'b01010100110111011110: color_data = 12'b111011101110;
20'b01010100110111011111: color_data = 12'b111011101110;
20'b01010100110111100000: color_data = 12'b111011101110;
20'b01010100110111100001: color_data = 12'b111011101110;
20'b01010100110111100010: color_data = 12'b111011101110;
20'b01010100110111100011: color_data = 12'b111011101110;
20'b01010100110111100100: color_data = 12'b111011101110;
20'b01010100110111100101: color_data = 12'b111011101110;
20'b01010100110111100110: color_data = 12'b111011101110;
20'b01010100110111100111: color_data = 12'b111011101110;
20'b01010101000010100001: color_data = 12'b111011101110;
20'b01010101000010100010: color_data = 12'b111011101110;
20'b01010101000010100011: color_data = 12'b111011101110;
20'b01010101000010100100: color_data = 12'b111011101110;
20'b01010101000010100101: color_data = 12'b111011101110;
20'b01010101000010100110: color_data = 12'b111011101110;
20'b01010101000010100111: color_data = 12'b111011101110;
20'b01010101000010101000: color_data = 12'b111011101110;
20'b01010101000010101001: color_data = 12'b111011101110;
20'b01010101000010101010: color_data = 12'b111011101110;
20'b01010101000010101100: color_data = 12'b111011101110;
20'b01010101000010101101: color_data = 12'b111011101110;
20'b01010101000010101110: color_data = 12'b111011101110;
20'b01010101000010101111: color_data = 12'b111011101110;
20'b01010101000010110000: color_data = 12'b111011101110;
20'b01010101000010110001: color_data = 12'b111011101110;
20'b01010101000010110010: color_data = 12'b111011101110;
20'b01010101000010110011: color_data = 12'b111011101110;
20'b01010101000010110100: color_data = 12'b111011101110;
20'b01010101000010110101: color_data = 12'b111011101110;
20'b01010101000010110111: color_data = 12'b111011101110;
20'b01010101000010111000: color_data = 12'b111011101110;
20'b01010101000010111001: color_data = 12'b111011101110;
20'b01010101000010111010: color_data = 12'b111011101110;
20'b01010101000010111011: color_data = 12'b111011101110;
20'b01010101000010111100: color_data = 12'b111011101110;
20'b01010101000010111101: color_data = 12'b111011101110;
20'b01010101000010111110: color_data = 12'b111011101110;
20'b01010101000010111111: color_data = 12'b111011101110;
20'b01010101000011000000: color_data = 12'b111011101110;
20'b01010101000011000010: color_data = 12'b111011101110;
20'b01010101000011000011: color_data = 12'b111011101110;
20'b01010101000011000100: color_data = 12'b111011101110;
20'b01010101000011000101: color_data = 12'b111011101110;
20'b01010101000011000110: color_data = 12'b111011101110;
20'b01010101000011000111: color_data = 12'b111011101110;
20'b01010101000011001000: color_data = 12'b111011101110;
20'b01010101000011001001: color_data = 12'b111011101110;
20'b01010101000011001010: color_data = 12'b111011101110;
20'b01010101000011001011: color_data = 12'b111011101110;
20'b01010101000011001101: color_data = 12'b111011101110;
20'b01010101000011001110: color_data = 12'b111011101110;
20'b01010101000011001111: color_data = 12'b111011101110;
20'b01010101000011010000: color_data = 12'b111011101110;
20'b01010101000011010001: color_data = 12'b111011101110;
20'b01010101000011010010: color_data = 12'b111011101110;
20'b01010101000011010011: color_data = 12'b111011101110;
20'b01010101000011010100: color_data = 12'b111011101110;
20'b01010101000011010101: color_data = 12'b111011101110;
20'b01010101000011010110: color_data = 12'b111011101110;
20'b01010101000100000011: color_data = 12'b111011101110;
20'b01010101000100000100: color_data = 12'b111011101110;
20'b01010101000100000101: color_data = 12'b111011101110;
20'b01010101000100000110: color_data = 12'b111011101110;
20'b01010101000100000111: color_data = 12'b111011101110;
20'b01010101000100001000: color_data = 12'b111011101110;
20'b01010101000100001001: color_data = 12'b111011101110;
20'b01010101000100001010: color_data = 12'b111011101110;
20'b01010101000100001011: color_data = 12'b111011101110;
20'b01010101000100001100: color_data = 12'b111011101110;
20'b01010101000100001110: color_data = 12'b111011101110;
20'b01010101000100001111: color_data = 12'b111011101110;
20'b01010101000100010000: color_data = 12'b111011101110;
20'b01010101000100010001: color_data = 12'b111011101110;
20'b01010101000100010010: color_data = 12'b111011101110;
20'b01010101000100010011: color_data = 12'b111011101110;
20'b01010101000100010100: color_data = 12'b111011101110;
20'b01010101000100010101: color_data = 12'b111011101110;
20'b01010101000100010110: color_data = 12'b111011101110;
20'b01010101000100010111: color_data = 12'b111011101110;
20'b01010101000100011001: color_data = 12'b111011101110;
20'b01010101000100011010: color_data = 12'b111011101110;
20'b01010101000100011011: color_data = 12'b111011101110;
20'b01010101000100011100: color_data = 12'b111011101110;
20'b01010101000100011101: color_data = 12'b111011101110;
20'b01010101000100011110: color_data = 12'b111011101110;
20'b01010101000100011111: color_data = 12'b111011101110;
20'b01010101000100100000: color_data = 12'b111011101110;
20'b01010101000100100001: color_data = 12'b111011101110;
20'b01010101000100100010: color_data = 12'b111011101110;
20'b01010101000101000100: color_data = 12'b111011101110;
20'b01010101000101000101: color_data = 12'b111011101110;
20'b01010101000101000110: color_data = 12'b111011101110;
20'b01010101000101000111: color_data = 12'b111011101110;
20'b01010101000101001000: color_data = 12'b111011101110;
20'b01010101000101001001: color_data = 12'b111011101110;
20'b01010101000101001010: color_data = 12'b111011101110;
20'b01010101000101001011: color_data = 12'b111011101110;
20'b01010101000101001100: color_data = 12'b111011101110;
20'b01010101000101001101: color_data = 12'b111011101110;
20'b01010101000101001111: color_data = 12'b111011101110;
20'b01010101000101010000: color_data = 12'b111011101110;
20'b01010101000101010001: color_data = 12'b111011101110;
20'b01010101000101010010: color_data = 12'b111011101110;
20'b01010101000101010011: color_data = 12'b111011101110;
20'b01010101000101010100: color_data = 12'b111011101110;
20'b01010101000101010101: color_data = 12'b111011101110;
20'b01010101000101010110: color_data = 12'b111011101110;
20'b01010101000101010111: color_data = 12'b111011101110;
20'b01010101000101011000: color_data = 12'b111011101110;
20'b01010101000101011010: color_data = 12'b111011101110;
20'b01010101000101011011: color_data = 12'b111011101110;
20'b01010101000101011100: color_data = 12'b111011101110;
20'b01010101000101011101: color_data = 12'b111011101110;
20'b01010101000101011110: color_data = 12'b111011101110;
20'b01010101000101011111: color_data = 12'b111011101110;
20'b01010101000101100000: color_data = 12'b111011101110;
20'b01010101000101100001: color_data = 12'b111011101110;
20'b01010101000101100010: color_data = 12'b111011101110;
20'b01010101000101100011: color_data = 12'b111011101110;
20'b01010101000101100101: color_data = 12'b111011101110;
20'b01010101000101100110: color_data = 12'b111011101110;
20'b01010101000101100111: color_data = 12'b111011101110;
20'b01010101000101101000: color_data = 12'b111011101110;
20'b01010101000101101001: color_data = 12'b111011101110;
20'b01010101000101101010: color_data = 12'b111011101110;
20'b01010101000101101011: color_data = 12'b111011101110;
20'b01010101000101101100: color_data = 12'b111011101110;
20'b01010101000101101101: color_data = 12'b111011101110;
20'b01010101000101101110: color_data = 12'b111011101110;
20'b01010101000101110000: color_data = 12'b111011101110;
20'b01010101000101110001: color_data = 12'b111011101110;
20'b01010101000101110010: color_data = 12'b111011101110;
20'b01010101000101110011: color_data = 12'b111011101110;
20'b01010101000101110100: color_data = 12'b111011101110;
20'b01010101000101110101: color_data = 12'b111011101110;
20'b01010101000101110110: color_data = 12'b111011101110;
20'b01010101000101110111: color_data = 12'b111011101110;
20'b01010101000101111000: color_data = 12'b111011101110;
20'b01010101000101111001: color_data = 12'b111011101110;
20'b01010101000101111011: color_data = 12'b111011101110;
20'b01010101000101111100: color_data = 12'b111011101110;
20'b01010101000101111101: color_data = 12'b111011101110;
20'b01010101000101111110: color_data = 12'b111011101110;
20'b01010101000101111111: color_data = 12'b111011101110;
20'b01010101000110000000: color_data = 12'b111011101110;
20'b01010101000110000001: color_data = 12'b111011101110;
20'b01010101000110000010: color_data = 12'b111011101110;
20'b01010101000110000011: color_data = 12'b111011101110;
20'b01010101000110000100: color_data = 12'b111011101110;
20'b01010101000110000110: color_data = 12'b111011101110;
20'b01010101000110000111: color_data = 12'b111011101110;
20'b01010101000110001000: color_data = 12'b111011101110;
20'b01010101000110001001: color_data = 12'b111011101110;
20'b01010101000110001010: color_data = 12'b111011101110;
20'b01010101000110001011: color_data = 12'b111011101110;
20'b01010101000110001100: color_data = 12'b111011101110;
20'b01010101000110001101: color_data = 12'b111011101110;
20'b01010101000110001110: color_data = 12'b111011101110;
20'b01010101000110001111: color_data = 12'b111011101110;
20'b01010101000110011100: color_data = 12'b111011101110;
20'b01010101000110011101: color_data = 12'b111011101110;
20'b01010101000110011110: color_data = 12'b111011101110;
20'b01010101000110011111: color_data = 12'b111011101110;
20'b01010101000110100000: color_data = 12'b111011101110;
20'b01010101000110100001: color_data = 12'b111011101110;
20'b01010101000110100010: color_data = 12'b111011101110;
20'b01010101000110100011: color_data = 12'b111011101110;
20'b01010101000110100100: color_data = 12'b111011101110;
20'b01010101000110100101: color_data = 12'b111011101110;
20'b01010101000110100111: color_data = 12'b111011101110;
20'b01010101000110101000: color_data = 12'b111011101110;
20'b01010101000110101001: color_data = 12'b111011101110;
20'b01010101000110101010: color_data = 12'b111011101110;
20'b01010101000110101011: color_data = 12'b111011101110;
20'b01010101000110101100: color_data = 12'b111011101110;
20'b01010101000110101101: color_data = 12'b111011101110;
20'b01010101000110101110: color_data = 12'b111011101110;
20'b01010101000110101111: color_data = 12'b111011101110;
20'b01010101000110110000: color_data = 12'b111011101110;
20'b01010101000111010011: color_data = 12'b111011101110;
20'b01010101000111010100: color_data = 12'b111011101110;
20'b01010101000111010101: color_data = 12'b111011101110;
20'b01010101000111010110: color_data = 12'b111011101110;
20'b01010101000111010111: color_data = 12'b111011101110;
20'b01010101000111011000: color_data = 12'b111011101110;
20'b01010101000111011001: color_data = 12'b111011101110;
20'b01010101000111011010: color_data = 12'b111011101110;
20'b01010101000111011011: color_data = 12'b111011101110;
20'b01010101000111011100: color_data = 12'b111011101110;
20'b01010101000111011110: color_data = 12'b111011101110;
20'b01010101000111011111: color_data = 12'b111011101110;
20'b01010101000111100000: color_data = 12'b111011101110;
20'b01010101000111100001: color_data = 12'b111011101110;
20'b01010101000111100010: color_data = 12'b111011101110;
20'b01010101000111100011: color_data = 12'b111011101110;
20'b01010101000111100100: color_data = 12'b111011101110;
20'b01010101000111100101: color_data = 12'b111011101110;
20'b01010101000111100110: color_data = 12'b111011101110;
20'b01010101000111100111: color_data = 12'b111011101110;
20'b01010101010010100001: color_data = 12'b111011101110;
20'b01010101010010100010: color_data = 12'b111011101110;
20'b01010101010010100011: color_data = 12'b111011101110;
20'b01010101010010100100: color_data = 12'b111011101110;
20'b01010101010010100101: color_data = 12'b111011101110;
20'b01010101010010100110: color_data = 12'b111011101110;
20'b01010101010010100111: color_data = 12'b111011101110;
20'b01010101010010101000: color_data = 12'b111011101110;
20'b01010101010010101001: color_data = 12'b111011101110;
20'b01010101010010101010: color_data = 12'b111011101110;
20'b01010101010010101100: color_data = 12'b111011101110;
20'b01010101010010101101: color_data = 12'b111011101110;
20'b01010101010010101110: color_data = 12'b111011101110;
20'b01010101010010101111: color_data = 12'b111011101110;
20'b01010101010010110000: color_data = 12'b111011101110;
20'b01010101010010110001: color_data = 12'b111011101110;
20'b01010101010010110010: color_data = 12'b111011101110;
20'b01010101010010110011: color_data = 12'b111011101110;
20'b01010101010010110100: color_data = 12'b111011101110;
20'b01010101010010110101: color_data = 12'b111011101110;
20'b01010101010010110111: color_data = 12'b111011101110;
20'b01010101010010111000: color_data = 12'b111011101110;
20'b01010101010010111001: color_data = 12'b111011101110;
20'b01010101010010111010: color_data = 12'b111011101110;
20'b01010101010010111011: color_data = 12'b111011101110;
20'b01010101010010111100: color_data = 12'b111011101110;
20'b01010101010010111101: color_data = 12'b111011101110;
20'b01010101010010111110: color_data = 12'b111011101110;
20'b01010101010010111111: color_data = 12'b111011101110;
20'b01010101010011000000: color_data = 12'b111011101110;
20'b01010101010011000010: color_data = 12'b111011101110;
20'b01010101010011000011: color_data = 12'b111011101110;
20'b01010101010011000100: color_data = 12'b111011101110;
20'b01010101010011000101: color_data = 12'b111011101110;
20'b01010101010011000110: color_data = 12'b111011101110;
20'b01010101010011000111: color_data = 12'b111011101110;
20'b01010101010011001000: color_data = 12'b111011101110;
20'b01010101010011001001: color_data = 12'b111011101110;
20'b01010101010011001010: color_data = 12'b111011101110;
20'b01010101010011001011: color_data = 12'b111011101110;
20'b01010101010011001101: color_data = 12'b111011101110;
20'b01010101010011001110: color_data = 12'b111011101110;
20'b01010101010011001111: color_data = 12'b111011101110;
20'b01010101010011010000: color_data = 12'b111011101110;
20'b01010101010011010001: color_data = 12'b111011101110;
20'b01010101010011010010: color_data = 12'b111011101110;
20'b01010101010011010011: color_data = 12'b111011101110;
20'b01010101010011010100: color_data = 12'b111011101110;
20'b01010101010011010101: color_data = 12'b111011101110;
20'b01010101010011010110: color_data = 12'b111011101110;
20'b01010101010100000011: color_data = 12'b111011101110;
20'b01010101010100000100: color_data = 12'b111011101110;
20'b01010101010100000101: color_data = 12'b111011101110;
20'b01010101010100000110: color_data = 12'b111011101110;
20'b01010101010100000111: color_data = 12'b111011101110;
20'b01010101010100001000: color_data = 12'b111011101110;
20'b01010101010100001001: color_data = 12'b111011101110;
20'b01010101010100001010: color_data = 12'b111011101110;
20'b01010101010100001011: color_data = 12'b111011101110;
20'b01010101010100001100: color_data = 12'b111011101110;
20'b01010101010100001110: color_data = 12'b111011101110;
20'b01010101010100001111: color_data = 12'b111011101110;
20'b01010101010100010000: color_data = 12'b111011101110;
20'b01010101010100010001: color_data = 12'b111011101110;
20'b01010101010100010010: color_data = 12'b111011101110;
20'b01010101010100010011: color_data = 12'b111011101110;
20'b01010101010100010100: color_data = 12'b111011101110;
20'b01010101010100010101: color_data = 12'b111011101110;
20'b01010101010100010110: color_data = 12'b111011101110;
20'b01010101010100010111: color_data = 12'b111011101110;
20'b01010101010100011001: color_data = 12'b111011101110;
20'b01010101010100011010: color_data = 12'b111011101110;
20'b01010101010100011011: color_data = 12'b111011101110;
20'b01010101010100011100: color_data = 12'b111011101110;
20'b01010101010100011101: color_data = 12'b111011101110;
20'b01010101010100011110: color_data = 12'b111011101110;
20'b01010101010100011111: color_data = 12'b111011101110;
20'b01010101010100100000: color_data = 12'b111011101110;
20'b01010101010100100001: color_data = 12'b111011101110;
20'b01010101010100100010: color_data = 12'b111011101110;
20'b01010101010101000100: color_data = 12'b111011101110;
20'b01010101010101000101: color_data = 12'b111011101110;
20'b01010101010101000110: color_data = 12'b111011101110;
20'b01010101010101000111: color_data = 12'b111011101110;
20'b01010101010101001000: color_data = 12'b111011101110;
20'b01010101010101001001: color_data = 12'b111011101110;
20'b01010101010101001010: color_data = 12'b111011101110;
20'b01010101010101001011: color_data = 12'b111011101110;
20'b01010101010101001100: color_data = 12'b111011101110;
20'b01010101010101001101: color_data = 12'b111011101110;
20'b01010101010101001111: color_data = 12'b111011101110;
20'b01010101010101010000: color_data = 12'b111011101110;
20'b01010101010101010001: color_data = 12'b111011101110;
20'b01010101010101010010: color_data = 12'b111011101110;
20'b01010101010101010011: color_data = 12'b111011101110;
20'b01010101010101010100: color_data = 12'b111011101110;
20'b01010101010101010101: color_data = 12'b111011101110;
20'b01010101010101010110: color_data = 12'b111011101110;
20'b01010101010101010111: color_data = 12'b111011101110;
20'b01010101010101011000: color_data = 12'b111011101110;
20'b01010101010101011010: color_data = 12'b111011101110;
20'b01010101010101011011: color_data = 12'b111011101110;
20'b01010101010101011100: color_data = 12'b111011101110;
20'b01010101010101011101: color_data = 12'b111011101110;
20'b01010101010101011110: color_data = 12'b111011101110;
20'b01010101010101011111: color_data = 12'b111011101110;
20'b01010101010101100000: color_data = 12'b111011101110;
20'b01010101010101100001: color_data = 12'b111011101110;
20'b01010101010101100010: color_data = 12'b111011101110;
20'b01010101010101100011: color_data = 12'b111011101110;
20'b01010101010101100101: color_data = 12'b111011101110;
20'b01010101010101100110: color_data = 12'b111011101110;
20'b01010101010101100111: color_data = 12'b111011101110;
20'b01010101010101101000: color_data = 12'b111011101110;
20'b01010101010101101001: color_data = 12'b111011101110;
20'b01010101010101101010: color_data = 12'b111011101110;
20'b01010101010101101011: color_data = 12'b111011101110;
20'b01010101010101101100: color_data = 12'b111011101110;
20'b01010101010101101101: color_data = 12'b111011101110;
20'b01010101010101101110: color_data = 12'b111011101110;
20'b01010101010101110000: color_data = 12'b111011101110;
20'b01010101010101110001: color_data = 12'b111011101110;
20'b01010101010101110010: color_data = 12'b111011101110;
20'b01010101010101110011: color_data = 12'b111011101110;
20'b01010101010101110100: color_data = 12'b111011101110;
20'b01010101010101110101: color_data = 12'b111011101110;
20'b01010101010101110110: color_data = 12'b111011101110;
20'b01010101010101110111: color_data = 12'b111011101110;
20'b01010101010101111000: color_data = 12'b111011101110;
20'b01010101010101111001: color_data = 12'b111011101110;
20'b01010101010101111011: color_data = 12'b111011101110;
20'b01010101010101111100: color_data = 12'b111011101110;
20'b01010101010101111101: color_data = 12'b111011101110;
20'b01010101010101111110: color_data = 12'b111011101110;
20'b01010101010101111111: color_data = 12'b111011101110;
20'b01010101010110000000: color_data = 12'b111011101110;
20'b01010101010110000001: color_data = 12'b111011101110;
20'b01010101010110000010: color_data = 12'b111011101110;
20'b01010101010110000011: color_data = 12'b111011101110;
20'b01010101010110000100: color_data = 12'b111011101110;
20'b01010101010110000110: color_data = 12'b111011101110;
20'b01010101010110000111: color_data = 12'b111011101110;
20'b01010101010110001000: color_data = 12'b111011101110;
20'b01010101010110001001: color_data = 12'b111011101110;
20'b01010101010110001010: color_data = 12'b111011101110;
20'b01010101010110001011: color_data = 12'b111011101110;
20'b01010101010110001100: color_data = 12'b111011101110;
20'b01010101010110001101: color_data = 12'b111011101110;
20'b01010101010110001110: color_data = 12'b111011101110;
20'b01010101010110001111: color_data = 12'b111011101110;
20'b01010101010110011100: color_data = 12'b111011101110;
20'b01010101010110011101: color_data = 12'b111011101110;
20'b01010101010110011110: color_data = 12'b111011101110;
20'b01010101010110011111: color_data = 12'b111011101110;
20'b01010101010110100000: color_data = 12'b111011101110;
20'b01010101010110100001: color_data = 12'b111011101110;
20'b01010101010110100010: color_data = 12'b111011101110;
20'b01010101010110100011: color_data = 12'b111011101110;
20'b01010101010110100100: color_data = 12'b111011101110;
20'b01010101010110100101: color_data = 12'b111011101110;
20'b01010101010110100111: color_data = 12'b111011101110;
20'b01010101010110101000: color_data = 12'b111011101110;
20'b01010101010110101001: color_data = 12'b111011101110;
20'b01010101010110101010: color_data = 12'b111011101110;
20'b01010101010110101011: color_data = 12'b111011101110;
20'b01010101010110101100: color_data = 12'b111011101110;
20'b01010101010110101101: color_data = 12'b111011101110;
20'b01010101010110101110: color_data = 12'b111011101110;
20'b01010101010110101111: color_data = 12'b111011101110;
20'b01010101010110110000: color_data = 12'b111011101110;
20'b01010101010111010011: color_data = 12'b111011101110;
20'b01010101010111010100: color_data = 12'b111011101110;
20'b01010101010111010101: color_data = 12'b111011101110;
20'b01010101010111010110: color_data = 12'b111011101110;
20'b01010101010111010111: color_data = 12'b111011101110;
20'b01010101010111011000: color_data = 12'b111011101110;
20'b01010101010111011001: color_data = 12'b111011101110;
20'b01010101010111011010: color_data = 12'b111011101110;
20'b01010101010111011011: color_data = 12'b111011101110;
20'b01010101010111011100: color_data = 12'b111011101110;
20'b01010101010111011110: color_data = 12'b111011101110;
20'b01010101010111011111: color_data = 12'b111011101110;
20'b01010101010111100000: color_data = 12'b111011101110;
20'b01010101010111100001: color_data = 12'b111011101110;
20'b01010101010111100010: color_data = 12'b111011101110;
20'b01010101010111100011: color_data = 12'b111011101110;
20'b01010101010111100100: color_data = 12'b111011101110;
20'b01010101010111100101: color_data = 12'b111011101110;
20'b01010101010111100110: color_data = 12'b111011101110;
20'b01010101010111100111: color_data = 12'b111011101110;
20'b01010101100010100001: color_data = 12'b111011101110;
20'b01010101100010100010: color_data = 12'b111011101110;
20'b01010101100010100011: color_data = 12'b111011101110;
20'b01010101100010100100: color_data = 12'b111011101110;
20'b01010101100010100101: color_data = 12'b111011101110;
20'b01010101100010100110: color_data = 12'b111011101110;
20'b01010101100010100111: color_data = 12'b111011101110;
20'b01010101100010101000: color_data = 12'b111011101110;
20'b01010101100010101001: color_data = 12'b111011101110;
20'b01010101100010101010: color_data = 12'b111011101110;
20'b01010101100010101100: color_data = 12'b111011101110;
20'b01010101100010101101: color_data = 12'b111011101110;
20'b01010101100010101110: color_data = 12'b111011101110;
20'b01010101100010101111: color_data = 12'b111011101110;
20'b01010101100010110000: color_data = 12'b111011101110;
20'b01010101100010110001: color_data = 12'b111011101110;
20'b01010101100010110010: color_data = 12'b111011101110;
20'b01010101100010110011: color_data = 12'b111011101110;
20'b01010101100010110100: color_data = 12'b111011101110;
20'b01010101100010110101: color_data = 12'b111011101110;
20'b01010101100010110111: color_data = 12'b111011101110;
20'b01010101100010111000: color_data = 12'b111011101110;
20'b01010101100010111001: color_data = 12'b111011101110;
20'b01010101100010111010: color_data = 12'b111011101110;
20'b01010101100010111011: color_data = 12'b111011101110;
20'b01010101100010111100: color_data = 12'b111011101110;
20'b01010101100010111101: color_data = 12'b111011101110;
20'b01010101100010111110: color_data = 12'b111011101110;
20'b01010101100010111111: color_data = 12'b111011101110;
20'b01010101100011000000: color_data = 12'b111011101110;
20'b01010101100011000010: color_data = 12'b111011101110;
20'b01010101100011000011: color_data = 12'b111011101110;
20'b01010101100011000100: color_data = 12'b111011101110;
20'b01010101100011000101: color_data = 12'b111011101110;
20'b01010101100011000110: color_data = 12'b111011101110;
20'b01010101100011000111: color_data = 12'b111011101110;
20'b01010101100011001000: color_data = 12'b111011101110;
20'b01010101100011001001: color_data = 12'b111011101110;
20'b01010101100011001010: color_data = 12'b111011101110;
20'b01010101100011001011: color_data = 12'b111011101110;
20'b01010101100011001101: color_data = 12'b111011101110;
20'b01010101100011001110: color_data = 12'b111011101110;
20'b01010101100011001111: color_data = 12'b111011101110;
20'b01010101100011010000: color_data = 12'b111011101110;
20'b01010101100011010001: color_data = 12'b111011101110;
20'b01010101100011010010: color_data = 12'b111011101110;
20'b01010101100011010011: color_data = 12'b111011101110;
20'b01010101100011010100: color_data = 12'b111011101110;
20'b01010101100011010101: color_data = 12'b111011101110;
20'b01010101100011010110: color_data = 12'b111011101110;
20'b01010101100100000011: color_data = 12'b111011101110;
20'b01010101100100000100: color_data = 12'b111011101110;
20'b01010101100100000101: color_data = 12'b111011101110;
20'b01010101100100000110: color_data = 12'b111011101110;
20'b01010101100100000111: color_data = 12'b111011101110;
20'b01010101100100001000: color_data = 12'b111011101110;
20'b01010101100100001001: color_data = 12'b111011101110;
20'b01010101100100001010: color_data = 12'b111011101110;
20'b01010101100100001011: color_data = 12'b111011101110;
20'b01010101100100001100: color_data = 12'b111011101110;
20'b01010101100100001110: color_data = 12'b111011101110;
20'b01010101100100001111: color_data = 12'b111011101110;
20'b01010101100100010000: color_data = 12'b111011101110;
20'b01010101100100010001: color_data = 12'b111011101110;
20'b01010101100100010010: color_data = 12'b111011101110;
20'b01010101100100010011: color_data = 12'b111011101110;
20'b01010101100100010100: color_data = 12'b111011101110;
20'b01010101100100010101: color_data = 12'b111011101110;
20'b01010101100100010110: color_data = 12'b111011101110;
20'b01010101100100010111: color_data = 12'b111011101110;
20'b01010101100100011001: color_data = 12'b111011101110;
20'b01010101100100011010: color_data = 12'b111011101110;
20'b01010101100100011011: color_data = 12'b111011101110;
20'b01010101100100011100: color_data = 12'b111011101110;
20'b01010101100100011101: color_data = 12'b111011101110;
20'b01010101100100011110: color_data = 12'b111011101110;
20'b01010101100100011111: color_data = 12'b111011101110;
20'b01010101100100100000: color_data = 12'b111011101110;
20'b01010101100100100001: color_data = 12'b111011101110;
20'b01010101100100100010: color_data = 12'b111011101110;
20'b01010101100101000100: color_data = 12'b111011101110;
20'b01010101100101000101: color_data = 12'b111011101110;
20'b01010101100101000110: color_data = 12'b111011101110;
20'b01010101100101000111: color_data = 12'b111011101110;
20'b01010101100101001000: color_data = 12'b111011101110;
20'b01010101100101001001: color_data = 12'b111011101110;
20'b01010101100101001010: color_data = 12'b111011101110;
20'b01010101100101001011: color_data = 12'b111011101110;
20'b01010101100101001100: color_data = 12'b111011101110;
20'b01010101100101001101: color_data = 12'b111011101110;
20'b01010101100101001111: color_data = 12'b111011101110;
20'b01010101100101010000: color_data = 12'b111011101110;
20'b01010101100101010001: color_data = 12'b111011101110;
20'b01010101100101010010: color_data = 12'b111011101110;
20'b01010101100101010011: color_data = 12'b111011101110;
20'b01010101100101010100: color_data = 12'b111011101110;
20'b01010101100101010101: color_data = 12'b111011101110;
20'b01010101100101010110: color_data = 12'b111011101110;
20'b01010101100101010111: color_data = 12'b111011101110;
20'b01010101100101011000: color_data = 12'b111011101110;
20'b01010101100101011010: color_data = 12'b111011101110;
20'b01010101100101011011: color_data = 12'b111011101110;
20'b01010101100101011100: color_data = 12'b111011101110;
20'b01010101100101011101: color_data = 12'b111011101110;
20'b01010101100101011110: color_data = 12'b111011101110;
20'b01010101100101011111: color_data = 12'b111011101110;
20'b01010101100101100000: color_data = 12'b111011101110;
20'b01010101100101100001: color_data = 12'b111011101110;
20'b01010101100101100010: color_data = 12'b111011101110;
20'b01010101100101100011: color_data = 12'b111011101110;
20'b01010101100101100101: color_data = 12'b111011101110;
20'b01010101100101100110: color_data = 12'b111011101110;
20'b01010101100101100111: color_data = 12'b111011101110;
20'b01010101100101101000: color_data = 12'b111011101110;
20'b01010101100101101001: color_data = 12'b111011101110;
20'b01010101100101101010: color_data = 12'b111011101110;
20'b01010101100101101011: color_data = 12'b111011101110;
20'b01010101100101101100: color_data = 12'b111011101110;
20'b01010101100101101101: color_data = 12'b111011101110;
20'b01010101100101101110: color_data = 12'b111011101110;
20'b01010101100101110000: color_data = 12'b111011101110;
20'b01010101100101110001: color_data = 12'b111011101110;
20'b01010101100101110010: color_data = 12'b111011101110;
20'b01010101100101110011: color_data = 12'b111011101110;
20'b01010101100101110100: color_data = 12'b111011101110;
20'b01010101100101110101: color_data = 12'b111011101110;
20'b01010101100101110110: color_data = 12'b111011101110;
20'b01010101100101110111: color_data = 12'b111011101110;
20'b01010101100101111000: color_data = 12'b111011101110;
20'b01010101100101111001: color_data = 12'b111011101110;
20'b01010101100101111011: color_data = 12'b111011101110;
20'b01010101100101111100: color_data = 12'b111011101110;
20'b01010101100101111101: color_data = 12'b111011101110;
20'b01010101100101111110: color_data = 12'b111011101110;
20'b01010101100101111111: color_data = 12'b111011101110;
20'b01010101100110000000: color_data = 12'b111011101110;
20'b01010101100110000001: color_data = 12'b111011101110;
20'b01010101100110000010: color_data = 12'b111011101110;
20'b01010101100110000011: color_data = 12'b111011101110;
20'b01010101100110000100: color_data = 12'b111011101110;
20'b01010101100110000110: color_data = 12'b111011101110;
20'b01010101100110000111: color_data = 12'b111011101110;
20'b01010101100110001000: color_data = 12'b111011101110;
20'b01010101100110001001: color_data = 12'b111011101110;
20'b01010101100110001010: color_data = 12'b111011101110;
20'b01010101100110001011: color_data = 12'b111011101110;
20'b01010101100110001100: color_data = 12'b111011101110;
20'b01010101100110001101: color_data = 12'b111011101110;
20'b01010101100110001110: color_data = 12'b111011101110;
20'b01010101100110001111: color_data = 12'b111011101110;
20'b01010101100110011100: color_data = 12'b111011101110;
20'b01010101100110011101: color_data = 12'b111011101110;
20'b01010101100110011110: color_data = 12'b111011101110;
20'b01010101100110011111: color_data = 12'b111011101110;
20'b01010101100110100000: color_data = 12'b111011101110;
20'b01010101100110100001: color_data = 12'b111011101110;
20'b01010101100110100010: color_data = 12'b111011101110;
20'b01010101100110100011: color_data = 12'b111011101110;
20'b01010101100110100100: color_data = 12'b111011101110;
20'b01010101100110100101: color_data = 12'b111011101110;
20'b01010101100110100111: color_data = 12'b111011101110;
20'b01010101100110101000: color_data = 12'b111011101110;
20'b01010101100110101001: color_data = 12'b111011101110;
20'b01010101100110101010: color_data = 12'b111011101110;
20'b01010101100110101011: color_data = 12'b111011101110;
20'b01010101100110101100: color_data = 12'b111011101110;
20'b01010101100110101101: color_data = 12'b111011101110;
20'b01010101100110101110: color_data = 12'b111011101110;
20'b01010101100110101111: color_data = 12'b111011101110;
20'b01010101100110110000: color_data = 12'b111011101110;
20'b01010101100111010011: color_data = 12'b111011101110;
20'b01010101100111010100: color_data = 12'b111011101110;
20'b01010101100111010101: color_data = 12'b111011101110;
20'b01010101100111010110: color_data = 12'b111011101110;
20'b01010101100111010111: color_data = 12'b111011101110;
20'b01010101100111011000: color_data = 12'b111011101110;
20'b01010101100111011001: color_data = 12'b111011101110;
20'b01010101100111011010: color_data = 12'b111011101110;
20'b01010101100111011011: color_data = 12'b111011101110;
20'b01010101100111011100: color_data = 12'b111011101110;
20'b01010101100111011110: color_data = 12'b111011101110;
20'b01010101100111011111: color_data = 12'b111011101110;
20'b01010101100111100000: color_data = 12'b111011101110;
20'b01010101100111100001: color_data = 12'b111011101110;
20'b01010101100111100010: color_data = 12'b111011101110;
20'b01010101100111100011: color_data = 12'b111011101110;
20'b01010101100111100100: color_data = 12'b111011101110;
20'b01010101100111100101: color_data = 12'b111011101110;
20'b01010101100111100110: color_data = 12'b111011101110;
20'b01010101100111100111: color_data = 12'b111011101110;
default: color_data = 12'b0;


	endcase
	end
endmodule